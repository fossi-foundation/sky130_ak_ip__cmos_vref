magic
tech sky130A
magscale 1 2
timestamp 1713056482
<< pwell >>
rect -1288 -3227 1288 3227
<< psubdiff >>
rect -1252 3157 -1156 3191
rect 1156 3157 1252 3191
rect -1252 3095 -1218 3157
rect 1218 3095 1252 3157
rect -1252 -3157 -1218 -3095
rect 1218 -3157 1252 -3095
rect -1252 -3191 -1156 -3157
rect 1156 -3191 1252 -3157
<< psubdiffcont >>
rect -1156 3157 1156 3191
rect -1252 -3095 -1218 3095
rect 1218 -3095 1252 3095
rect -1156 -3191 1156 -3157
<< xpolycontact >>
rect -1122 2629 -984 3061
rect -1122 -3061 -984 -2629
rect -888 2629 -750 3061
rect -888 -3061 -750 -2629
rect -654 2629 -516 3061
rect -654 -3061 -516 -2629
rect -420 2629 -282 3061
rect -420 -3061 -282 -2629
rect -186 2629 -48 3061
rect -186 -3061 -48 -2629
rect 48 2629 186 3061
rect 48 -3061 186 -2629
rect 282 2629 420 3061
rect 282 -3061 420 -2629
rect 516 2629 654 3061
rect 516 -3061 654 -2629
rect 750 2629 888 3061
rect 750 -3061 888 -2629
rect 984 2629 1122 3061
rect 984 -3061 1122 -2629
<< xpolyres >>
rect -1122 -2629 -984 2629
rect -888 -2629 -750 2629
rect -654 -2629 -516 2629
rect -420 -2629 -282 2629
rect -186 -2629 -48 2629
rect 48 -2629 186 2629
rect 282 -2629 420 2629
rect 516 -2629 654 2629
rect 750 -2629 888 2629
rect 984 -2629 1122 2629
<< locali >>
rect -1252 3157 -1156 3191
rect 1156 3157 1252 3191
rect -1252 3095 -1218 3157
rect 1218 3095 1252 3157
rect -1252 -3157 -1218 -3095
rect 1218 -3157 1252 -3095
rect -1252 -3191 -1156 -3157
rect 1156 -3191 1252 -3157
<< viali >>
rect -1106 2646 -1000 3043
rect -872 2646 -766 3043
rect -638 2646 -532 3043
rect -404 2646 -298 3043
rect -170 2646 -64 3043
rect 64 2646 170 3043
rect 298 2646 404 3043
rect 532 2646 638 3043
rect 766 2646 872 3043
rect 1000 2646 1106 3043
rect -1106 -3043 -1000 -2646
rect -872 -3043 -766 -2646
rect -638 -3043 -532 -2646
rect -404 -3043 -298 -2646
rect -170 -3043 -64 -2646
rect 64 -3043 170 -2646
rect 298 -3043 404 -2646
rect 532 -3043 638 -2646
rect 766 -3043 872 -2646
rect 1000 -3043 1106 -2646
<< metal1 >>
rect -1112 3043 -994 3055
rect -1112 2646 -1106 3043
rect -1000 2646 -994 3043
rect -1112 2634 -994 2646
rect -878 3043 -760 3055
rect -878 2646 -872 3043
rect -766 2646 -760 3043
rect -878 2634 -760 2646
rect -644 3043 -526 3055
rect -644 2646 -638 3043
rect -532 2646 -526 3043
rect -644 2634 -526 2646
rect -410 3043 -292 3055
rect -410 2646 -404 3043
rect -298 2646 -292 3043
rect -410 2634 -292 2646
rect -176 3043 -58 3055
rect -176 2646 -170 3043
rect -64 2646 -58 3043
rect -176 2634 -58 2646
rect 58 3043 176 3055
rect 58 2646 64 3043
rect 170 2646 176 3043
rect 58 2634 176 2646
rect 292 3043 410 3055
rect 292 2646 298 3043
rect 404 2646 410 3043
rect 292 2634 410 2646
rect 526 3043 644 3055
rect 526 2646 532 3043
rect 638 2646 644 3043
rect 526 2634 644 2646
rect 760 3043 878 3055
rect 760 2646 766 3043
rect 872 2646 878 3043
rect 760 2634 878 2646
rect 994 3043 1112 3055
rect 994 2646 1000 3043
rect 1106 2646 1112 3043
rect 994 2634 1112 2646
rect -1112 -2646 -994 -2634
rect -1112 -3043 -1106 -2646
rect -1000 -3043 -994 -2646
rect -1112 -3055 -994 -3043
rect -878 -2646 -760 -2634
rect -878 -3043 -872 -2646
rect -766 -3043 -760 -2646
rect -878 -3055 -760 -3043
rect -644 -2646 -526 -2634
rect -644 -3043 -638 -2646
rect -532 -3043 -526 -2646
rect -644 -3055 -526 -3043
rect -410 -2646 -292 -2634
rect -410 -3043 -404 -2646
rect -298 -3043 -292 -2646
rect -410 -3055 -292 -3043
rect -176 -2646 -58 -2634
rect -176 -3043 -170 -2646
rect -64 -3043 -58 -2646
rect -176 -3055 -58 -3043
rect 58 -2646 176 -2634
rect 58 -3043 64 -2646
rect 170 -3043 176 -2646
rect 58 -3055 176 -3043
rect 292 -2646 410 -2634
rect 292 -3043 298 -2646
rect 404 -3043 410 -2646
rect 292 -3055 410 -3043
rect 526 -2646 644 -2634
rect 526 -3043 532 -2646
rect 638 -3043 644 -2646
rect 526 -3055 644 -3043
rect 760 -2646 878 -2634
rect 760 -3043 766 -2646
rect 872 -3043 878 -2646
rect 760 -3055 878 -3043
rect 994 -2646 1112 -2634
rect 994 -3043 1000 -2646
rect 1106 -3043 1112 -2646
rect 994 -3055 1112 -3043
<< properties >>
string FIXED_BBOX -1235 -3174 1235 3174
string gencell sky130_fd_pr__res_xhigh_po_0p69
string library sky130
string parameters w 0.690 l 26.45 m 1 nx 10 wmin 0.690 lmin 0.50 rho 2000 val 77.212k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.690 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
