magic
tech sky130A
magscale 1 2
timestamp 1713045697
<< error_p >>
rect -1011 263 1031 274
rect -984 254 1031 263
rect -1112 240 1112 254
rect -1160 164 -1126 219
rect -1046 200 -1012 204
rect 1012 200 1046 204
rect -1080 172 -1062 178
rect -1058 172 -1006 200
rect 984 182 1058 200
rect -994 178 1058 182
rect -996 172 1058 178
rect 1062 172 1080 178
rect -1084 138 -1006 172
rect -1000 138 1084 172
rect 1126 164 1160 219
rect -1080 132 -1062 138
rect -1058 104 -1006 138
rect -996 132 996 138
rect -994 128 994 132
rect 1006 104 1058 138
rect 1062 132 1080 138
rect -1058 100 -1036 104
rect -1022 100 -1012 104
rect 1012 100 1022 104
rect 1036 100 1058 104
rect -1058 -104 -1036 -100
rect -1022 -104 -1012 -100
rect 984 -104 1022 -100
rect 1036 -104 1058 -100
rect -1080 -138 -1062 -132
rect -1058 -138 -1006 -104
rect 984 -128 1058 -104
rect -994 -132 1058 -128
rect -996 -138 1058 -132
rect 1062 -138 1080 -132
rect -1084 -141 -1006 -138
rect -1126 -164 -1006 -141
rect -1160 -172 -1006 -164
rect -1000 -172 1084 -138
rect 1160 -164 1207 -141
rect 1126 -172 1207 -164
rect -1160 -199 -1126 -172
rect -1080 -178 -1062 -172
rect -1058 -186 -1006 -172
rect -996 -178 996 -172
rect -994 -182 994 -178
rect 1006 -186 1058 -172
rect 1062 -178 1080 -172
rect -1058 -200 -1000 -186
rect 1000 -200 1058 -186
rect 1126 -199 1160 -172
rect -1046 -204 -1012 -200
rect 1012 -204 1046 -200
rect -984 -238 984 -206
rect -1011 -250 1011 -240
rect -1011 -251 -984 -250
rect 984 -251 1011 -250
rect -1000 -263 1000 -258
rect -1011 -274 1011 -263
<< pwell >>
rect -1196 310 1196 410
rect -5312 -310 5312 310
rect -1196 -410 1196 -310
<< nmos >>
rect -5116 -100 -3116 100
rect -3058 -100 -1058 100
rect -1000 172 1000 200
rect -1000 138 -984 172
rect 984 138 1000 172
rect -1000 -138 1000 138
rect -1000 -172 -984 -138
rect 984 -172 1000 -138
rect -1000 -200 1000 -172
rect 1058 -100 3058 100
rect 3116 -100 5116 100
<< ndiff >>
rect -1058 188 -1000 200
rect -5174 88 -5116 100
rect -5174 -88 -5162 88
rect -5128 -88 -5116 88
rect -5174 -100 -5116 -88
rect -3116 88 -3058 100
rect -3116 -88 -3104 88
rect -3070 -88 -3058 88
rect -3116 -100 -3058 -88
rect -1058 -188 -1046 188
rect -1012 -188 -1000 188
rect 1000 188 1058 200
rect -1058 -200 -1000 -188
rect 1000 -188 1012 188
rect 1046 -188 1058 188
rect 3058 88 3116 100
rect 3058 -88 3070 88
rect 3104 -88 3116 88
rect 3058 -100 3116 -88
rect 5116 88 5174 100
rect 5116 -88 5128 88
rect 5162 -88 5174 88
rect 5116 -100 5174 -88
rect 1000 -200 1058 -188
<< ndiffc >>
rect -5162 -88 -5128 88
rect -3104 -88 -3070 88
rect -1046 -188 -1012 188
rect 1012 -188 1046 188
rect 3070 -88 3104 88
rect 5128 -88 5162 88
<< psubdiff >>
rect -1160 340 -1064 374
rect 1064 340 1160 374
rect -1160 278 -1126 340
rect 1126 278 1160 340
rect -5276 240 -5180 274
rect 5180 240 5276 274
rect -5276 178 -5242 240
rect -5276 -240 -5242 -178
rect 5242 178 5276 240
rect 5242 -240 5276 -178
rect -5276 -274 -5180 -240
rect 5180 -274 5276 -240
rect -1160 -340 -1126 -278
rect 1126 -340 1160 -278
rect -1160 -374 -1064 -340
rect 1064 -374 1160 -340
<< psubdiffcont >>
rect -1064 340 1064 374
rect -1160 274 -1126 278
rect 1126 274 1160 278
rect -5180 240 5180 274
rect -1160 188 -1126 240
rect -5276 -178 -5242 178
rect 1126 188 1160 240
rect -1160 -240 -1126 -188
rect 5242 -178 5276 178
rect 1126 -240 1160 -188
rect -5180 -274 5180 -240
rect -1160 -278 -1126 -274
rect 1126 -278 1160 -274
rect -1064 -374 1064 -340
<< poly >>
rect -1000 274 1000 288
rect -1000 238 -984 240
rect 984 238 1000 240
rect -1000 200 1000 238
rect -5116 172 -3116 188
rect -5116 138 -5100 172
rect -3132 138 -3116 172
rect -5116 100 -3116 138
rect -3058 172 -1058 188
rect -3058 138 -3042 172
rect -1074 138 -1058 172
rect -3058 100 -1058 138
rect -5116 -138 -3116 -100
rect -5116 -172 -5100 -138
rect -3132 -172 -3116 -138
rect -5116 -188 -3116 -172
rect -3058 -138 -1058 -100
rect -3058 -172 -3042 -138
rect -1074 -172 -1058 -138
rect -3058 -188 -1058 -172
rect 1058 172 3058 188
rect 1058 138 1074 172
rect 3042 138 3058 172
rect 1058 100 3058 138
rect 3116 172 5116 188
rect 3116 138 3132 172
rect 5100 138 5116 172
rect 3116 100 5116 138
rect 1058 -138 3058 -100
rect 1058 -172 1074 -138
rect 3042 -172 3058 -138
rect 1058 -188 3058 -172
rect 3116 -138 5116 -100
rect 3116 -172 3132 -138
rect 5100 -172 5116 -138
rect 3116 -188 5116 -172
rect -1000 -238 1000 -200
rect -1000 -240 -984 -238
rect 984 -240 1000 -238
rect -1000 -288 1000 -274
<< polycont >>
rect -984 238 984 240
rect -5100 138 -3132 172
rect -3042 138 -1074 172
rect -5100 -172 -3132 -138
rect -3042 -172 -1074 -138
rect -984 138 984 172
rect -984 -172 984 -138
rect 1074 138 3042 172
rect 3132 138 5100 172
rect 1074 -172 3042 -138
rect 3132 -172 5100 -138
rect -984 -240 984 -238
<< locali >>
rect -1160 340 -1064 374
rect 1064 340 1160 374
rect -1160 278 -1126 340
rect 1126 278 1160 340
rect -5276 240 -5180 274
rect 5180 240 5276 274
rect -5276 178 -5242 240
rect -1000 238 -984 240
rect 984 238 1000 240
rect -1160 172 -1126 188
rect -1046 188 -1012 204
rect -5116 138 -5100 172
rect -3132 138 -3116 172
rect -3058 138 -3042 172
rect -1074 138 -1058 172
rect -5162 88 -5128 104
rect -5162 -104 -5128 -88
rect -3104 88 -3070 104
rect -3104 -104 -3070 -88
rect -1160 -138 -1126 138
rect -5116 -172 -5100 -138
rect -3132 -172 -3116 -138
rect -3058 -172 -3042 -138
rect -1074 -172 -1058 -138
rect -5276 -240 -5242 -178
rect -1160 -188 -1126 -172
rect 1012 188 1046 204
rect -1000 138 -984 172
rect 984 138 1000 172
rect -1000 -172 -984 -138
rect 984 -172 1000 -138
rect -1046 -204 -1012 -188
rect 1126 172 1160 188
rect 5242 178 5276 240
rect 1058 138 1074 172
rect 3042 138 3058 172
rect 3116 138 3132 172
rect 5100 138 5116 172
rect 1126 -138 1160 138
rect 3070 88 3104 104
rect 3070 -104 3104 -88
rect 5128 88 5162 104
rect 5128 -104 5162 -88
rect 1058 -172 1074 -138
rect 3042 -172 3058 -138
rect 3116 -172 3132 -138
rect 5100 -172 5116 -138
rect 1012 -204 1046 -188
rect 1126 -188 1160 -172
rect -1000 -240 -984 -238
rect 984 -240 1000 -238
rect 5242 -240 5276 -178
rect -5276 -274 -5180 -240
rect 5180 -274 5276 -240
rect -1160 -340 -1126 -278
rect 1126 -340 1160 -278
rect -1160 -374 -1064 -340
rect 1064 -374 1160 -340
<< viali >>
rect -984 240 984 272
rect -984 238 984 240
rect -5100 138 -3132 172
rect -3042 138 -1074 172
rect -5162 -88 -5128 88
rect -3104 -88 -3070 88
rect -5100 -172 -3132 -138
rect -3042 -172 -1074 -138
rect -1046 -188 -1012 188
rect -984 138 984 172
rect -984 -172 984 -138
rect 1012 -188 1046 188
rect 1074 138 3042 172
rect 3132 138 5100 172
rect 3070 -88 3104 88
rect 5128 -88 5162 88
rect 1074 -172 3042 -138
rect 3132 -172 5100 -138
rect -984 -240 984 -238
rect -984 -272 984 -240
<< metal1 >>
rect -996 272 996 278
rect -996 238 -984 272
rect 984 238 996 272
rect -996 232 996 238
rect -1052 188 -1006 200
rect -5112 172 -3120 178
rect -5112 138 -5100 172
rect -3132 138 -3120 172
rect -5112 132 -3120 138
rect -3054 172 -1062 178
rect -3054 138 -3042 172
rect -1074 138 -1062 172
rect -3054 132 -1062 138
rect -5168 88 -5122 100
rect -5168 -88 -5162 88
rect -5128 -88 -5122 88
rect -5168 -100 -5122 -88
rect -3110 88 -3064 100
rect -3110 -88 -3104 88
rect -3070 -88 -3064 88
rect -3110 -100 -3064 -88
rect -5112 -138 -3120 -132
rect -5112 -172 -5100 -138
rect -3132 -172 -3120 -138
rect -5112 -178 -3120 -172
rect -3054 -138 -1062 -132
rect -3054 -172 -3042 -138
rect -1074 -172 -1062 -138
rect -3054 -178 -1062 -172
rect -1052 -188 -1046 188
rect -1012 -188 -1006 188
rect 1006 188 1052 200
rect -996 172 996 178
rect -996 138 -984 172
rect 984 138 996 172
rect -996 132 996 138
rect -996 -138 996 -132
rect -996 -172 -984 -138
rect 984 -172 996 -138
rect -996 -178 996 -172
rect -1052 -200 -1006 -188
rect 1006 -188 1012 188
rect 1046 -188 1052 188
rect 1062 172 3054 178
rect 1062 138 1074 172
rect 3042 138 3054 172
rect 1062 132 3054 138
rect 3120 172 5112 178
rect 3120 138 3132 172
rect 5100 138 5112 172
rect 3120 132 5112 138
rect 3064 88 3110 100
rect 3064 -88 3070 88
rect 3104 -88 3110 88
rect 3064 -100 3110 -88
rect 5122 88 5168 100
rect 5122 -88 5128 88
rect 5162 -88 5168 88
rect 5122 -100 5168 -88
rect 1062 -138 3054 -132
rect 1062 -172 1074 -138
rect 3042 -172 3054 -138
rect 1062 -178 3054 -172
rect 3120 -138 5112 -132
rect 3120 -172 3132 -138
rect 5100 -172 5112 -138
rect 3120 -178 5112 -172
rect 1006 -200 1052 -188
rect -996 -238 996 -232
rect -996 -272 -984 -238
rect 984 -272 996 -238
rect -996 -278 996 -272
<< properties >>
string FIXED_BBOX -5259 -257 5259 257
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.0 l 10.0 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
