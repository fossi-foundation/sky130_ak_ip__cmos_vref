magic
tech sky130A
timestamp 1713212409
<< pwell >>
rect -348 -355 348 355
<< nmos >>
rect -250 -250 250 250
<< ndiff >>
rect -279 244 -250 250
rect -279 -244 -273 244
rect -256 -244 -250 244
rect -279 -250 -250 -244
rect 250 244 279 250
rect 250 -244 256 244
rect 273 -244 279 244
rect 250 -250 279 -244
<< ndiffc >>
rect -273 -244 -256 244
rect 256 -244 273 244
<< psubdiff >>
rect -330 320 -282 337
rect 282 320 330 337
rect -330 289 -313 320
rect 313 289 330 320
rect -330 -320 -313 -289
rect 313 -320 330 -289
rect -330 -337 -282 -320
rect 282 -337 330 -320
<< psubdiffcont >>
rect -282 320 282 337
rect -330 -289 -313 289
rect 313 -289 330 289
rect -282 -337 282 -320
<< poly >>
rect -250 286 250 294
rect -250 269 -242 286
rect 242 269 250 286
rect -250 250 250 269
rect -250 -269 250 -250
rect -250 -286 -242 -269
rect 242 -286 250 -269
rect -250 -294 250 -286
<< polycont >>
rect -242 269 242 286
rect -242 -286 242 -269
<< locali >>
rect -330 320 -282 337
rect 282 320 330 337
rect -330 289 -313 320
rect 313 289 330 320
rect -250 269 -242 286
rect 242 269 250 286
rect -273 244 -256 252
rect -273 -252 -256 -244
rect 256 244 273 252
rect 256 -252 273 -244
rect -250 -286 -242 -269
rect 242 -286 250 -269
rect -330 -320 -313 -289
rect 313 -320 330 -289
rect -330 -337 -282 -320
rect 282 -337 330 -320
<< viali >>
rect -242 269 242 286
rect -273 -244 -256 244
rect 256 -244 273 244
rect -242 -286 242 -269
<< metal1 >>
rect -248 286 248 289
rect -248 269 -242 286
rect 242 269 248 286
rect -248 266 248 269
rect -276 244 -253 250
rect -276 -244 -273 244
rect -256 -244 -253 244
rect -276 -250 -253 -244
rect 253 244 276 250
rect 253 -244 256 244
rect 273 -244 276 244
rect 253 -250 276 -244
rect -248 -269 248 -266
rect -248 -286 -242 -269
rect 242 -286 248 -269
rect -248 -289 248 -286
<< properties >>
string FIXED_BBOX -321 -328 321 328
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 5 l 5.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
