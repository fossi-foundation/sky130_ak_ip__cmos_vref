magic
tech sky130A
magscale 1 2
timestamp 1716240972
<< error_s >>
rect 14489 -5908 14515 -5903
rect 13794 -6200 13800 -6194
rect 13800 -6206 13806 -6200
rect 19600 -11708 19606 -11702
rect 19794 -11708 19800 -11702
rect 19594 -11714 19600 -11708
rect 19800 -11714 19806 -11708
rect 10112 -17190 10115 -16908
rect 10140 -17218 10143 -16880
<< metal1 >>
rect 9219 -400 14900 -200
rect 9068 -4238 9132 -450
rect 9219 -2449 11719 -2443
rect 9219 -2501 9225 -2449
rect 11713 -2501 11719 -2449
rect 9219 -2507 11719 -2501
rect 9068 -4482 9074 -4238
rect 9126 -4482 9132 -4238
rect 9068 -4488 9132 -4482
rect 11805 -4250 11869 -450
rect 11955 -2449 14455 -2443
rect 11955 -2501 11961 -2449
rect 14449 -2501 14455 -2449
rect 11955 -2507 14455 -2501
rect 11805 -4494 11811 -4250
rect 11863 -4494 11869 -4250
rect 14542 -4238 14606 -450
rect 14542 -4482 14548 -4238
rect 14600 -4482 14606 -4238
rect 14542 -4488 14606 -4482
rect 14700 -3400 14900 -400
rect 15000 -781 15200 -200
rect 15300 -400 15500 -200
rect 15391 -691 15460 -400
rect 15391 -734 15400 -691
rect 15394 -743 15400 -734
rect 15452 -734 15460 -691
rect 15452 -743 15458 -734
rect 15394 -749 15458 -743
rect 15000 -981 15344 -781
rect 15216 -2781 15344 -981
rect 15500 -1300 15700 -781
rect 15494 -1500 15700 -1300
rect 15500 -1700 16000 -1500
rect 15393 -2820 15459 -2812
rect 15393 -2872 15400 -2820
rect 15452 -2872 15459 -2820
rect 15393 -2878 15459 -2872
rect 15500 -3400 15700 -1700
rect 14700 -3600 15700 -3400
rect 11805 -4500 11869 -4494
rect 9219 -4620 11719 -4556
rect 11955 -4620 14455 -4556
rect 14700 -4620 14900 -3600
rect 15000 -3700 15200 -3694
rect 15200 -3900 15400 -3700
rect 15000 -3906 15400 -3900
rect 15200 -4280 15400 -3906
rect 15180 -4300 15420 -4280
rect 15180 -4500 15200 -4300
rect 15400 -4500 15420 -4300
rect 15180 -4520 15420 -4500
rect 9220 -4820 14900 -4620
rect 13780 -5000 14020 -4980
rect 15200 -5000 15400 -4520
rect 13780 -5148 13800 -5000
rect 9300 -5200 13800 -5148
rect 14000 -5200 15400 -5000
rect 9300 -5212 14020 -5200
rect 13780 -5220 14020 -5212
rect 8999 -5790 9290 -5289
rect 13302 -5300 13450 -5286
rect 13302 -5500 15200 -5300
rect 15400 -5500 15406 -5300
rect 9000 -8900 9200 -5790
rect 13302 -5794 13450 -5500
rect 9300 -5932 13864 -5868
rect 14206 -5898 14414 -5500
rect 13800 -6000 13864 -5932
rect 14487 -5969 14489 -5903
rect 14131 -6000 14489 -5969
rect 14000 -6200 14489 -6000
rect 12614 -6500 12700 -6300
rect 12900 -6500 13400 -6300
rect 13600 -6500 13623 -6300
rect 12700 -6504 13623 -6500
rect 13500 -6700 13700 -6694
rect 12500 -6900 13500 -6700
rect 12500 -8400 12700 -6900
rect 13500 -8400 13700 -6900
rect 14131 -7900 14489 -6200
rect 15500 -6300 15700 -3600
rect 15800 -4000 16000 -1800
rect 15800 -4206 16000 -4200
rect 15800 -4300 16000 -4294
rect 15800 -4506 16000 -4500
rect 14594 -6500 14600 -6300
rect 14800 -6500 15700 -6300
rect 14880 -7900 15120 -7880
rect 14131 -8100 14900 -7900
rect 15100 -8100 15120 -7900
rect 14880 -8120 15120 -8100
rect 14300 -8400 15200 -8200
rect 15400 -8400 15406 -8200
rect 12700 -8600 13600 -8500
rect 14300 -8600 14500 -8400
rect 12700 -8800 14500 -8600
rect 14580 -8600 14820 -8580
rect 15500 -8600 15700 -6500
rect 14580 -8800 14600 -8600
rect 14800 -8800 15700 -8600
rect 15800 -5300 16000 -5294
rect 15800 -8700 16000 -5500
rect 14580 -8820 14820 -8800
rect 15800 -8900 19000 -8700
rect 19200 -8900 19206 -8700
rect 9000 -9100 14300 -8900
rect 14500 -9100 15700 -8900
rect 9172 -9456 13000 -9338
rect 13205 -9456 14800 -9338
rect 12900 -9572 13000 -9456
rect 9172 -9924 9593 -9572
rect 12900 -9690 13626 -9572
rect 13205 -9924 14500 -9806
rect 9172 -10656 9593 -10304
rect 13297 -10422 14200 -10304
rect 9172 -11124 9593 -10772
rect 13297 -10890 13718 -10538
rect 14000 -10700 14200 -10422
rect 14300 -10400 14500 -9924
rect 14600 -10100 14800 -9456
rect 15500 -9500 15700 -9100
rect 19600 -9482 19800 -8679
rect 19578 -9500 19816 -9482
rect 15500 -9700 19600 -9500
rect 19800 -9700 19816 -9500
rect 19578 -9721 19816 -9700
rect 15194 -10000 15200 -9800
rect 15400 -10000 18700 -9800
rect 18900 -10000 18906 -9800
rect 18994 -10000 19000 -9800
rect 19200 -10000 21500 -9800
rect 14600 -10300 20500 -10100
rect 20700 -10300 21500 -10100
rect 17880 -10400 18120 -10380
rect 14300 -10600 17900 -10400
rect 18100 -10600 21500 -10400
rect 17880 -10620 18120 -10600
rect 14000 -10900 21500 -10700
rect 13297 -11124 14200 -11006
rect 14000 -11464 14200 -11124
rect 15800 -11400 16000 -10900
rect 9172 -11816 9593 -11464
rect 13351 -11582 15400 -11464
rect 17894 -11500 17900 -11300
rect 18100 -11500 18106 -11300
rect 9172 -12284 9593 -11932
rect 13351 -12050 13772 -11698
rect 14280 -11700 14520 -11680
rect 14280 -11900 14300 -11700
rect 14500 -11900 14520 -11700
rect 14280 -11920 14520 -11900
rect 14580 -11700 14820 -11680
rect 14580 -11900 14600 -11700
rect 14800 -11900 14820 -11700
rect 14580 -11920 14820 -11900
rect 14880 -11700 15120 -11680
rect 14880 -11900 14900 -11700
rect 15100 -11900 15120 -11700
rect 14880 -11920 15120 -11900
rect 9172 -12752 9593 -12400
rect 13351 -12518 13772 -12166
rect 9172 -13220 9593 -12868
rect 13351 -12986 13772 -12634
rect 9172 -13688 9593 -13336
rect 13351 -13454 13772 -13102
rect 9172 -14156 9593 -13804
rect 13351 -13922 13772 -13570
rect 9172 -14624 9593 -14272
rect 13351 -14390 13772 -14038
rect 11400 -14506 11600 -14500
rect 11400 -14624 13772 -14506
rect 9000 -15900 9200 -15700
rect 11400 -15900 11600 -14624
rect 14300 -14900 14500 -11920
rect 11900 -15100 14500 -14900
rect 11900 -15900 12100 -15100
rect 14600 -16608 14800 -11920
rect 14900 -16308 15100 -11920
rect 15200 -16008 15400 -11582
rect 18700 -11708 18900 -11702
rect 20480 -11708 20720 -11680
rect 20480 -11908 20500 -11708
rect 20700 -11908 20720 -11708
rect 18700 -11914 18900 -11908
rect 20480 -11920 20720 -11908
rect 15200 -16208 15700 -16008
rect 14900 -16508 15700 -16308
rect 14600 -16808 15700 -16608
rect 9000 -17600 9200 -17400
rect 9000 -17900 9200 -17700
rect 9000 -19500 9200 -19300
rect 14600 -19500 14800 -19300
rect 15200 -19500 15400 -19300
<< via1 >>
rect 9225 -2501 11713 -2449
rect 9074 -4482 9126 -4238
rect 11961 -2501 14449 -2449
rect 11811 -4494 11863 -4250
rect 14548 -4482 14600 -4238
rect 15400 -743 15452 -691
rect 15400 -2872 15452 -2820
rect 15000 -3900 15200 -3700
rect 15200 -4500 15400 -4300
rect 13800 -5200 14000 -5000
rect 15200 -5500 15400 -5300
rect 13800 -6200 14000 -6000
rect 12700 -6500 12900 -6300
rect 13400 -6500 13600 -6300
rect 13500 -6900 13700 -6700
rect 15800 -4200 16000 -4000
rect 15800 -4500 16000 -4300
rect 14600 -6500 14800 -6300
rect 14900 -8100 15100 -7900
rect 15200 -8400 15400 -8200
rect 14600 -8800 14800 -8600
rect 15800 -5500 16000 -5300
rect 19000 -8900 19200 -8700
rect 14300 -9100 14500 -8900
rect 19600 -9700 19800 -9500
rect 15200 -10000 15400 -9800
rect 18700 -10000 18900 -9800
rect 19000 -10000 19200 -9800
rect 20500 -10300 20700 -10100
rect 17900 -10600 18100 -10400
rect 17900 -11500 18100 -11300
rect 14300 -11900 14500 -11700
rect 14600 -11900 14800 -11700
rect 14900 -11900 15100 -11700
rect 18700 -11908 18900 -11708
rect 19600 -11908 19800 -11708
rect 20500 -11908 20700 -11708
<< metal2 >>
rect 15394 -691 15804 -685
rect 15394 -743 15400 -691
rect 15452 -743 15804 -691
rect 15394 -749 15804 -743
rect 9219 -2449 15200 -2411
rect 9219 -2501 9225 -2449
rect 11713 -2501 11961 -2449
rect 14449 -2501 15200 -2449
rect 9219 -2539 15200 -2501
rect 15000 -3700 15200 -2539
rect 15740 -2813 15804 -749
rect 15394 -2820 15804 -2813
rect 15394 -2872 15400 -2820
rect 15452 -2872 15804 -2820
rect 15394 -2877 15804 -2872
rect 14994 -3900 15000 -3700
rect 15200 -3900 15206 -3700
rect 14900 -4200 15800 -4000
rect 16000 -4200 16006 -4000
rect 9068 -4238 9132 -4232
rect 9068 -4482 9074 -4238
rect 9126 -4482 9132 -4238
rect 14542 -4238 14606 -4232
rect 9068 -4556 9132 -4482
rect 11805 -4250 11869 -4244
rect 11805 -4494 11811 -4250
rect 11863 -4494 11869 -4250
rect 11805 -4556 11869 -4494
rect 14542 -4482 14548 -4238
rect 14600 -4482 14606 -4238
rect 14542 -4556 14606 -4482
rect 14900 -4556 15100 -4200
rect 15180 -4300 15420 -4280
rect 15180 -4500 15200 -4300
rect 15400 -4500 15800 -4300
rect 16000 -4500 16006 -4300
rect 15180 -4520 15420 -4500
rect 9068 -4620 15100 -4556
rect 13780 -5000 14020 -4980
rect 13780 -5200 13800 -5000
rect 14000 -5200 14020 -5000
rect 13780 -5220 14020 -5200
rect 13800 -6000 14000 -5220
rect 13800 -6206 14000 -6200
rect 14600 -6300 14800 -6294
rect 12614 -6500 12700 -6300
rect 12900 -6500 13400 -6300
rect 13600 -6500 14600 -6300
rect 12700 -6504 13623 -6500
rect 13400 -6506 13600 -6504
rect 14600 -6506 14800 -6500
rect 14900 -6700 15100 -4620
rect 15200 -5300 15400 -5294
rect 15400 -5500 15800 -5300
rect 16000 -5500 16006 -5300
rect 15200 -5506 15400 -5500
rect 13494 -6900 13500 -6700
rect 13700 -6900 15100 -6700
rect 14880 -7900 15120 -7880
rect 14880 -8100 14900 -7900
rect 15100 -8100 15120 -7900
rect 14880 -8120 15120 -8100
rect 14580 -8600 14820 -8580
rect 14580 -8800 14600 -8600
rect 14800 -8800 14820 -8600
rect 14580 -8820 14820 -8800
rect 14300 -8900 14500 -8893
rect 14300 -11680 14500 -9100
rect 14600 -11680 14800 -8820
rect 14900 -11680 15100 -8120
rect 15200 -8200 15400 -8194
rect 15200 -9800 15400 -8400
rect 19000 -8700 19200 -8694
rect 15200 -10006 15400 -10000
rect 18700 -9800 18900 -9794
rect 17880 -10400 18120 -10380
rect 17880 -10600 17900 -10400
rect 18100 -10600 18120 -10400
rect 17880 -10620 18120 -10600
rect 17900 -11300 18100 -10620
rect 17900 -11506 18100 -11500
rect 14280 -11700 14520 -11680
rect 14280 -11900 14300 -11700
rect 14500 -11900 14520 -11700
rect 14280 -11920 14520 -11900
rect 14580 -11700 14820 -11680
rect 14580 -11900 14600 -11700
rect 14800 -11900 14820 -11700
rect 14580 -11920 14820 -11900
rect 14880 -11700 15120 -11680
rect 14880 -11900 14900 -11700
rect 15100 -11900 15120 -11700
rect 18700 -11708 18900 -10000
rect 19000 -9800 19200 -8900
rect 19578 -9500 19816 -9482
rect 19578 -9700 19600 -9500
rect 19800 -9700 19816 -9500
rect 19578 -9721 19816 -9700
rect 19000 -10006 19200 -10000
rect 19600 -11708 19800 -9721
rect 20500 -10100 20700 -10094
rect 20500 -11680 20700 -10300
rect 14880 -11920 15120 -11900
rect 18694 -11908 18700 -11708
rect 18900 -11908 18906 -11708
rect 20480 -11708 20720 -11680
rect 20480 -11908 20500 -11708
rect 20700 -11908 20720 -11708
rect 20480 -11920 20720 -11908
use sky130_fd_pr__res_xhigh_po_0p69_E9MCU4  R1
timestamp 1713140876
transform 0 1 11399 -1 0 -9631
box -469 -2399 469 2399
use sky130_fd_pr__res_xhigh_po_0p69_39QBTQ  R2
timestamp 1713056482
transform 0 1 16942 -1 0 -11365
box -235 -1442 235 1442
use sky130_fd_pr__res_xhigh_po_0p69_NB3ZKH  R3
timestamp 1713140876
transform 0 1 11445 -1 0 -10714
box -586 -2445 586 2445
use sky130_fd_pr__res_xhigh_po_0p69_GAZAU4  R4
timestamp 1713140876
transform 0 -1 11472 1 0 -13044
box -1756 -2472 1756 2472
use sbvfcm  x1
timestamp 1716240972
transform 1 0 10300 0 1 -5200
box 5700 -3700 11200 5000
use output_amp  x2
timestamp 1716240972
transform 1 0 10400 0 -1 -14608
box 5100 -2900 11120 4900
use trim_res  x3
timestamp 1713569381
transform 1 0 8300 0 1 -15600
box 700 -3900 5534 -100
use sky130_fd_pr__nfet_01v8_2333C8  XM1
timestamp 1713045697
transform 1 0 11296 0 1 -5540
box -2196 -460 2196 460
use sky130_fd_pr__nfet_01v8_QXBCRM  XM2
timestamp 1713051622
transform 0 -1 14310 1 0 -6904
box -1196 -310 1196 310
use sky130_fd_pr__pfet_01v8_6H4ZLK  XM3
timestamp 1716240972
transform 0 1 13119 -1 0 -7504
box -1196 -719 1196 719
use sky130_fd_pr__pfet_01v8_B3G3L7  XM9
timestamp 1713056482
transform 0 -1 11837 1 0 -2475
box -2225 -2837 2225 2837
use sky130_fd_pr__pfet_01v8_XPMKX6  XM20
timestamp 1713045697
transform 1 0 15426 0 1 -1781
box -226 -1219 226 1219
<< labels >>
flabel metal1 21300 -10300 21500 -10100 0 FreeSans 256 0 0 0 vbg
port 0 nsew
flabel metal1 21300 -10600 21500 -10400 0 FreeSans 256 0 0 0 vbgtg
port 7 nsew
flabel metal1 21300 -10900 21500 -10700 0 FreeSans 256 0 0 0 vbgsc
port 6 nsew
flabel metal1 9000 -9100 9200 -8900 0 FreeSans 256 0 0 0 avss
port 1 nsew
flabel metal1 21300 -10000 21500 -9800 0 FreeSans 256 0 0 0 vptat
port 13 nsew
flabel metal1 14600 -19500 14800 -19300 0 FreeSans 256 0 0 0 dvdd
port 3 nsew
flabel metal1 15200 -19500 15400 -19300 0 FreeSans 256 0 0 0 dvss
port 4 nsew
flabel metal1 9000 -19500 9200 -19300 0 FreeSans 256 0 0 0 trim3
port 8 nsew
flabel metal1 9000 -17900 9200 -17700 0 FreeSans 256 0 0 0 trim2
port 9 nsew
flabel metal1 9000 -17600 9200 -17400 0 FreeSans 256 0 0 0 trim1
port 10 nsew
flabel metal1 9000 -15900 9200 -15700 0 FreeSans 256 0 0 0 trim0
port 11 nsew
flabel metal1 15000 -400 15200 -200 0 FreeSans 256 0 0 0 avdd18
port 2 nsew
flabel metal1 15300 -400 15500 -200 0 FreeSans 256 0 0 0 ena
port 5 nsew
<< end >>
