magic
tech sky130A
magscale 1 2
timestamp 1716081120
<< nwell >>
rect -1225 -2219 1225 2219
<< pmos >>
rect -1029 -2000 -29 2000
rect 29 -2000 1029 2000
<< pdiff >>
rect -1087 1988 -1029 2000
rect -1087 -1988 -1075 1988
rect -1041 -1988 -1029 1988
rect -1087 -2000 -1029 -1988
rect -29 1988 29 2000
rect -29 -1988 -17 1988
rect 17 -1988 29 1988
rect -29 -2000 29 -1988
rect 1029 1988 1087 2000
rect 1029 -1988 1041 1988
rect 1075 -1988 1087 1988
rect 1029 -2000 1087 -1988
<< pdiffc >>
rect -1075 -1988 -1041 1988
rect -17 -1988 17 1988
rect 1041 -1988 1075 1988
<< nsubdiff >>
rect -1189 2149 -1093 2183
rect 1093 2149 1189 2183
rect -1189 2087 -1155 2149
rect 1155 2087 1189 2149
rect -1189 -2149 -1155 -2087
rect 1155 -2149 1189 -2087
rect -1189 -2183 -1093 -2149
rect 1093 -2183 1189 -2149
<< nsubdiffcont >>
rect -1093 2149 1093 2183
rect -1189 -2087 -1155 2087
rect 1155 -2087 1189 2087
rect -1093 -2183 1093 -2149
<< poly >>
rect -1029 2081 -29 2097
rect -1029 2047 -1013 2081
rect -45 2047 -29 2081
rect -1029 2000 -29 2047
rect 29 2081 1029 2097
rect 29 2047 45 2081
rect 1013 2047 1029 2081
rect 29 2000 1029 2047
rect -1029 -2047 -29 -2000
rect -1029 -2081 -1013 -2047
rect -45 -2081 -29 -2047
rect -1029 -2097 -29 -2081
rect 29 -2047 1029 -2000
rect 29 -2081 45 -2047
rect 1013 -2081 1029 -2047
rect 29 -2097 1029 -2081
<< polycont >>
rect -1013 2047 -45 2081
rect 45 2047 1013 2081
rect -1013 -2081 -45 -2047
rect 45 -2081 1013 -2047
<< locali >>
rect -1189 2149 -1093 2183
rect 1093 2149 1189 2183
rect -1189 2087 -1155 2149
rect 1155 2087 1189 2149
rect -1029 2047 -1013 2081
rect -45 2047 -29 2081
rect 29 2047 45 2081
rect 1013 2047 1029 2081
rect -1075 1988 -1041 2004
rect -1075 -2004 -1041 -1988
rect -17 1988 17 2004
rect -17 -2004 17 -1988
rect 1041 1988 1075 2004
rect 1041 -2004 1075 -1988
rect -1029 -2081 -1013 -2047
rect -45 -2081 -29 -2047
rect 29 -2081 45 -2047
rect 1013 -2081 1029 -2047
rect -1189 -2149 -1155 -2087
rect 1155 -2149 1189 -2087
rect -1189 -2183 -1093 -2149
rect 1093 -2183 1189 -2149
<< viali >>
rect -1013 2047 -45 2081
rect 45 2047 1013 2081
rect -1075 -1988 -1041 1988
rect -17 -1988 17 1988
rect 1041 -1988 1075 1988
rect -1013 -2081 -45 -2047
rect 45 -2081 1013 -2047
<< metal1 >>
rect -1025 2081 -33 2087
rect -1025 2047 -1013 2081
rect -45 2047 -33 2081
rect -1025 2041 -33 2047
rect 33 2081 1025 2087
rect 33 2047 45 2081
rect 1013 2047 1025 2081
rect 33 2041 1025 2047
rect -1081 1988 -1035 2000
rect -1081 -1988 -1075 1988
rect -1041 -1988 -1035 1988
rect -1081 -2000 -1035 -1988
rect -23 1988 23 2000
rect -23 -1988 -17 1988
rect 17 -1988 23 1988
rect -23 -2000 23 -1988
rect 1035 1988 1081 2000
rect 1035 -1988 1041 1988
rect 1075 -1988 1081 1988
rect 1035 -2000 1081 -1988
rect -1025 -2047 -33 -2041
rect -1025 -2081 -1013 -2047
rect -45 -2081 -33 -2047
rect -1025 -2087 -33 -2081
rect 33 -2047 1025 -2041
rect 33 -2081 45 -2047
rect 1013 -2081 1025 -2047
rect 33 -2087 1025 -2081
<< properties >>
string FIXED_BBOX -1172 -2166 1172 2166
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 20 l 5.0 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
