magic
tech sky130A
magscale 1 2
timestamp 1713051387
<< pwell >>
rect -201 -757 201 757
<< psubdiff >>
rect -165 687 -69 721
rect 69 687 165 721
rect -165 625 -131 687
rect 131 625 165 687
rect -165 -687 -131 -625
rect 131 -687 165 -625
rect -165 -721 -69 -687
rect 69 -721 165 -687
<< psubdiffcont >>
rect -69 687 69 721
rect -165 -625 -131 625
rect 131 -625 165 625
rect -69 -721 69 -687
<< xpolycontact >>
rect -35 159 35 591
rect -35 -591 35 -159
<< xpolyres >>
rect -35 -159 35 159
<< locali >>
rect -165 687 -69 721
rect 69 687 165 721
rect -165 625 -131 687
rect 131 625 165 687
rect -165 -687 -131 -625
rect 131 -687 165 -625
rect -165 -721 -69 -687
rect 69 -721 165 -687
<< viali >>
rect -19 176 19 573
rect -19 -573 19 -176
<< metal1 >>
rect -25 573 25 585
rect -25 176 -19 573
rect 19 176 25 573
rect -25 164 25 176
rect -25 -176 25 -164
rect -25 -573 -19 -176
rect 19 -573 25 -176
rect -25 -585 25 -573
<< properties >>
string FIXED_BBOX -148 -704 148 704
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 1.75 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 11.075k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
