magic
tech sky130A
magscale 1 2
timestamp 1713216111
<< error_p >>
rect 21300 -1594 21320 -1588
rect 21272 -1622 21292 -1616
rect 21274 -4500 21300 -4288
rect 21302 -4528 21328 -4260
rect 20500 -14708 20506 -14702
rect 20694 -14708 20700 -14702
rect 20494 -14714 20500 -14708
rect 20700 -14714 20706 -14708
rect 20494 -14908 20500 -14902
rect 20500 -14914 20506 -14908
<< error_s >>
rect 16372 -1594 16400 -1588
rect 16400 -1622 16428 -1616
rect 16294 -1894 16300 -1888
rect 16300 -1900 16306 -1894
rect 16300 -2094 16306 -2088
rect 16294 -2100 16300 -2094
rect 17300 -2194 17306 -2188
rect 17294 -2200 17300 -2194
rect 17294 -2394 17300 -2388
rect 17500 -2394 17506 -2388
rect 17300 -2400 17306 -2394
rect 17494 -2400 17500 -2394
rect 15597 -3328 15655 -3322
rect 15597 -3362 15609 -3328
rect 15597 -3368 15655 -3362
rect 17300 -3494 17306 -3488
rect 17294 -3500 17300 -3494
rect 17294 -3694 17300 -3688
rect 17300 -3700 17306 -3694
rect 18400 -4694 18420 -4688
rect 19272 -4694 19300 -4688
rect 18372 -4722 18392 -4716
rect 19300 -4722 19328 -4716
rect 19200 -5094 19206 -5088
rect 19394 -5094 19400 -5088
rect 19194 -5100 19200 -5094
rect 19400 -5100 19406 -5094
rect 19194 -5294 19200 -5288
rect 19400 -5294 19406 -5288
rect 19200 -5300 19206 -5294
rect 19394 -5300 19400 -5294
rect 19100 -5594 19106 -5588
rect 19294 -5594 19300 -5588
rect 19094 -5600 19100 -5594
rect 19300 -5600 19306 -5594
rect 19094 -5794 19100 -5788
rect 19100 -5800 19106 -5794
rect 19472 -6194 19500 -6188
rect 19500 -6222 19528 -6216
rect 18100 -6694 18106 -6688
rect 18294 -6694 18300 -6688
rect 18094 -6700 18100 -6694
rect 18300 -6700 18306 -6694
rect 18094 -6894 18100 -6888
rect 18300 -6894 18306 -6888
rect 18100 -6900 18106 -6894
rect 18294 -6900 18300 -6894
rect 18100 -7694 18106 -7688
rect 18294 -7694 18300 -7688
rect 18094 -7700 18100 -7694
rect 18300 -7700 18306 -7694
rect 18094 -7894 18100 -7888
rect 18300 -7894 18306 -7888
rect 18100 -7900 18106 -7894
rect 18294 -7900 18300 -7894
rect 14600 -8600 14606 -8594
rect 14594 -8606 14600 -8600
rect 14594 -8800 14600 -8794
rect 14600 -8806 14606 -8800
rect 19400 -9194 19406 -9188
rect 19594 -9194 19600 -9188
rect 19394 -9200 19400 -9194
rect 19600 -9200 19606 -9194
rect 19394 -9394 19400 -9388
rect 19600 -9394 19606 -9388
rect 19400 -9400 19406 -9394
rect 19594 -9400 19600 -9394
rect 19600 -9500 19606 -9494
rect 19794 -9500 19800 -9494
rect 19594 -9506 19600 -9500
rect 19800 -9506 19806 -9500
rect 17900 -10400 17906 -10394
rect 18094 -10400 18100 -10394
rect 17894 -10406 17900 -10400
rect 18100 -10406 18106 -10400
rect 14900 -11700 14906 -11694
rect 15094 -11700 15100 -11694
rect 14894 -11706 14900 -11700
rect 15100 -11706 15106 -11700
rect 19600 -11708 19606 -11702
rect 19794 -11708 19800 -11702
rect 19594 -11714 19600 -11708
rect 19800 -11714 19806 -11708
rect 14894 -11900 14900 -11894
rect 15100 -11900 15106 -11894
rect 14900 -11906 14906 -11900
rect 15094 -11906 15100 -11900
rect 19594 -11908 19600 -11902
rect 19800 -11908 19806 -11902
rect 19600 -11914 19606 -11908
rect 19794 -11914 19800 -11908
rect 17500 -12008 17506 -12002
rect 17694 -12008 17700 -12002
rect 17494 -12014 17500 -12008
rect 17700 -12014 17706 -12008
rect 17494 -12208 17500 -12202
rect 17700 -12208 17706 -12202
rect 17500 -12214 17506 -12208
rect 17694 -12214 17700 -12208
rect 19000 -13408 19006 -13402
rect 19194 -13408 19200 -13402
rect 18994 -13414 19000 -13408
rect 19200 -13414 19206 -13408
rect 18994 -13608 19000 -13602
rect 19200 -13608 19206 -13602
rect 19000 -13614 19006 -13608
rect 19194 -13614 19200 -13608
rect 10980 -16246 10986 -16240
rect 11174 -16246 11180 -16240
rect 10974 -16252 10980 -16246
rect 11180 -16252 11186 -16246
rect 10974 -16446 10980 -16440
rect 11180 -16446 11186 -16440
rect 10980 -16452 10986 -16446
rect 11174 -16452 11180 -16446
rect 14140 -16560 14146 -16554
rect 14334 -16560 14340 -16554
rect 14134 -16566 14140 -16560
rect 14340 -16566 14346 -16560
rect 13140 -16592 13146 -16586
rect 13146 -16598 13152 -16592
rect 14134 -16760 14140 -16755
rect 14340 -16760 14346 -16755
rect 14140 -16766 14146 -16760
rect 14334 -16766 14340 -16760
<< metal1 >>
rect 15200 -1900 15400 -700
rect 15500 -1200 15700 -700
rect 15200 -2100 15600 -1900
rect 15700 -2094 16100 -1894
rect 16000 -2394 16800 -2194
rect 15600 -3600 15800 -3594
rect 9000 -8500 9200 -8300
rect 15600 -8600 15800 -3800
rect 16000 -4900 16200 -2394
rect 16100 -5000 16300 -4994
rect 16100 -5206 16300 -5200
rect 9000 -8800 9200 -8600
rect 14800 -8800 15800 -8600
rect 9000 -9100 14300 -8900
rect 14500 -9100 16000 -8900
rect 13500 -9500 14800 -9300
rect 13500 -10000 14500 -9800
rect 13600 -10500 14200 -10300
rect 14000 -10700 14200 -10500
rect 14300 -10400 14500 -10000
rect 14600 -10100 14800 -9500
rect 15800 -9500 16000 -9100
rect 19700 -9500 19900 -9194
rect 15800 -9700 19600 -9500
rect 19800 -9700 19900 -9500
rect 17100 -10000 18700 -9800
rect 18900 -10000 18906 -9800
rect 20994 -10000 21000 -9800
rect 21200 -10000 21500 -9800
rect 14600 -10300 21500 -10100
rect 14300 -10600 17900 -10400
rect 18100 -10600 21500 -10400
rect 14000 -10900 21500 -10700
rect 15800 -11400 16000 -10900
rect 13600 -11600 15400 -11400
rect 17894 -11500 17900 -11300
rect 18100 -11500 18106 -11300
rect 14300 -11700 14500 -11694
rect 11640 -14700 13400 -14500
rect 11640 -15060 11840 -14700
rect 14300 -14860 14500 -11900
rect 11900 -15060 14500 -14860
rect 14600 -11700 14800 -11694
rect 9000 -15300 9200 -15100
rect 9000 -15600 9200 -15400
rect 14600 -16608 14800 -11900
rect 14900 -16308 15100 -11900
rect 15200 -16008 15400 -11600
rect 18700 -11708 18900 -11702
rect 18700 -11914 18900 -11908
rect 15200 -16208 15700 -16008
rect 14900 -16508 15700 -16308
rect 14600 -16808 15700 -16608
rect 9000 -19200 9200 -19000
rect 9000 -19500 9200 -19300
<< via1 >>
rect 16100 -2094 16300 -1894
rect 15600 -3800 15800 -3600
rect 16100 -5200 16300 -5000
rect 14600 -8800 14800 -8600
rect 14300 -9100 14500 -8900
rect 19400 -9394 19600 -9194
rect 19600 -9700 19800 -9500
rect 18700 -10000 18900 -9800
rect 21000 -10000 21200 -9800
rect 17900 -10600 18100 -10400
rect 17900 -11500 18100 -11300
rect 14300 -11900 14500 -11700
rect 14600 -11900 14800 -11700
rect 14900 -11900 15100 -11700
rect 18700 -11908 18900 -11708
rect 19600 -11908 19800 -11708
<< metal2 >>
rect 15700 -2094 16100 -1894
rect 15700 -3600 15900 -2094
rect 15594 -3800 15600 -3600
rect 15800 -3800 15900 -3600
rect 14900 -5200 16100 -5000
rect 16300 -5200 16306 -5000
rect 14600 -8600 14800 -8500
rect 14300 -8900 14500 -8893
rect 14300 -11700 14500 -9100
rect 14600 -11700 14800 -8800
rect 14900 -11700 15100 -5200
rect 19600 -9394 21200 -9194
rect 18700 -9800 18900 -9794
rect 17900 -11300 18100 -10600
rect 17900 -11506 18100 -11500
rect 14294 -11900 14300 -11700
rect 14500 -11900 14506 -11700
rect 14594 -11900 14600 -11700
rect 14800 -11900 14806 -11700
rect 18700 -11708 18900 -10000
rect 19600 -11708 19800 -9700
rect 21000 -9800 21200 -9394
rect 21000 -10006 21200 -10000
rect 18694 -11908 18700 -11708
rect 18900 -11908 18906 -11708
use sky130_fd_pr__res_xhigh_po_0p69_E9MCU4  R1
timestamp 1713140876
transform 0 1 11399 -1 0 -9631
box -469 -2399 469 2399
use sky130_fd_pr__res_xhigh_po_0p69_39QBTQ  R2
timestamp 1713056482
transform 0 1 16942 -1 0 -11365
box -235 -1442 235 1442
use sky130_fd_pr__res_xhigh_po_0p69_NB3ZKH  R3
timestamp 1713140876
transform 0 1 11445 -1 0 -10714
box -586 -2445 586 2445
use sky130_fd_pr__res_xhigh_po_0p69_GAZAU4  R4
timestamp 1713140876
transform 0 -1 11472 1 0 -13044
box -1756 -2472 1756 2472
use sbvfcm  x1
timestamp 1713214705
transform 1 0 10400 0 1 -5694
box 5700 -3706 11200 5500
use output_amp  x2
timestamp 1713128983
transform 1 0 10400 0 -1 -14608
box 5100 -2903 11100 4892
use trim_res  x3
timestamp 1713116496
transform 1 0 8480 0 1 -15320
box 720 -4180 5972 460
use sky130_fd_pr__nfet_01v8_2333C8  XM1
timestamp 1713045697
transform 1 0 11196 0 1 -5840
box -2196 -460 2196 460
use sky130_fd_pr__nfet_01v8_QXBCRM  XM2
timestamp 1713051622
transform 1 0 10196 0 1 -6690
box -1196 -310 1196 310
use sky130_fd_pr__pfet_01v8_6H4ZLK  XM3
timestamp 1713045697
transform 1 0 12696 0 1 -7081
box -1196 -719 1196 719
use sky130_fd_pr__pfet_01v8_B3G3L7  XM9
timestamp 1713056482
transform 0 -1 11937 1 0 -3075
box -2225 -2837 2225 2837
use sky130_fd_pr__pfet_01v8_XPMKX6  XM20
timestamp 1713045697
transform 1 0 15626 0 1 -2281
box -226 -1219 226 1219
<< labels >>
flabel metal1 21300 -10300 21500 -10100 0 FreeSans 256 0 0 0 vbg
port 0 nsew
flabel metal1 21300 -10600 21500 -10400 0 FreeSans 256 0 0 0 vbgtg
port 7 nsew
flabel metal1 21300 -10900 21500 -10700 0 FreeSans 256 0 0 0 vbgsc
port 6 nsew
flabel metal1 15500 -900 15700 -700 0 FreeSans 256 0 0 0 ena
port 5 nsew
flabel metal1 9000 -19500 9200 -19300 0 FreeSans 256 0 0 0 trim3
port 8 nsew
flabel metal1 9000 -19200 9200 -19000 0 FreeSans 256 0 0 0 trim2
port 9 nsew
flabel metal1 9000 -15600 9200 -15400 0 FreeSans 256 0 0 0 trim0
port 11 nsew
flabel metal1 9000 -15300 9200 -15100 0 FreeSans 256 0 0 0 trim1
port 10 nsew
flabel metal1 9000 -9100 9200 -8900 0 FreeSans 256 0 0 0 avss
port 1 nsew
flabel metal1 9000 -8800 9200 -8600 0 FreeSans 256 0 0 0 dvss
port 4 nsew
flabel metal1 9000 -8500 9200 -8300 0 FreeSans 256 0 0 0 dvdd
port 3 nsew
flabel metal1 21300 -10000 21500 -9800 0 FreeSans 256 0 0 0 vptat
port 13 nsew
flabel metal1 15200 -900 15400 -700 0 FreeSans 256 0 0 0 avdd18
port 2 nsew
<< end >>
