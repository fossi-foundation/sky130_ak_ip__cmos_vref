magic
tech sky130A
magscale 1 2
timestamp 1719454670
<< dnwell >>
rect 8800 -6220 21700 0
rect 11927 -9496 21700 -6220
rect 8800 -19700 21700 -9496
<< nwell >>
rect 8720 -1800 21780 80
rect 8720 -5955 9006 -1800
rect 8720 -5956 9331 -5955
rect 8720 -6300 12137 -5956
rect 8836 -7592 10984 -7553
rect 11792 -9308 12137 -6300
rect 8720 -9702 12137 -9308
rect 8720 -19494 9006 -9702
rect 21494 -15000 21780 -1800
rect 19000 -17100 21780 -15000
rect 15500 -19494 21780 -17100
rect 8720 -19780 21780 -19494
<< psubdiff >>
rect 8589 172 8649 206
rect 21861 172 21921 206
rect 8589 146 8623 172
rect 21887 146 21921 172
rect 8623 -6879 11516 -6869
rect 8623 -6908 8659 -6879
rect 8589 -6919 8659 -6908
rect 11414 -6919 11516 -6879
rect 8589 -6932 11516 -6919
rect 11453 -6968 11516 -6932
rect 8589 -7976 8623 -7946
rect 11453 -8916 11466 -6968
rect 11507 -8916 11516 -6968
rect 11453 -8950 11516 -8916
rect 8623 -8960 11516 -8950
rect 8623 -9000 8698 -8960
rect 11453 -9000 11516 -8960
rect 8623 -9013 11516 -9000
rect 8589 -19869 8623 -19843
rect 21887 -19869 21921 -19843
rect 8589 -19903 8649 -19869
rect 21861 -19903 21921 -19869
<< nsubdiff >>
rect 8757 23 21743 43
rect 8757 -11 8837 23
rect 21663 -11 21743 23
rect 8757 -31 21743 -11
rect 8757 -37 8831 -31
rect 8757 -6063 8777 -37
rect 8811 -6063 8831 -37
rect 8757 -6084 8831 -6063
rect 21669 -37 21743 -31
rect 8757 -6104 12054 -6084
rect 8757 -6138 8848 -6104
rect 11958 -6138 12054 -6104
rect 8757 -6158 12054 -6138
rect 11980 -6184 12054 -6158
rect 11980 -9527 11999 -6184
rect 12033 -9527 12054 -6184
rect 11980 -9546 12054 -9527
rect 8757 -9566 12054 -9546
rect 8757 -9600 8833 -9566
rect 11943 -9600 12054 -9566
rect 8757 -9620 12054 -9600
rect 8757 -9678 8831 -9620
rect 8757 -19663 8777 -9678
rect 8811 -19663 8831 -9678
rect 8757 -19669 8831 -19663
rect 21669 -19663 21689 -37
rect 21723 -19663 21743 -37
rect 21669 -19669 21743 -19663
rect 8757 -19689 21743 -19669
rect 8757 -19723 8837 -19689
rect 21663 -19723 21743 -19689
rect 8757 -19743 21743 -19723
<< psubdiffcont >>
rect 8649 172 21861 206
rect 8589 -6908 8623 146
rect 8659 -6919 11414 -6879
rect 8589 -19843 8623 -7976
rect 11466 -8916 11507 -6968
rect 8698 -9000 11453 -8960
rect 21887 -19843 21921 146
rect 8649 -19903 21861 -19869
<< nsubdiffcont >>
rect 8837 -11 21663 23
rect 8777 -6063 8811 -37
rect 8848 -6138 11958 -6104
rect 11999 -9527 12033 -6184
rect 8833 -9600 11943 -9566
rect 8777 -19663 8811 -9678
rect 21689 -19663 21723 -37
rect 8837 -19723 21663 -19689
<< locali >>
rect 8589 172 8649 206
rect 21861 172 21921 206
rect 8589 146 8715 172
rect 8623 132 8715 146
rect 21727 146 21921 172
rect 21727 139 21887 146
rect 21727 132 21860 139
rect 8623 108 21860 132
rect 8623 36 8678 108
rect 8651 -6093 8678 36
rect 8623 -6847 8678 -6093
rect 8737 34 21769 58
rect 8737 23 8869 34
rect 21623 23 21769 34
rect 8737 -11 8837 23
rect 21663 -11 21769 23
rect 8737 -18 8869 -11
rect 21623 -18 21769 -11
rect 8737 -37 21769 -18
rect 8737 -62 8777 -37
rect 8811 -47 21689 -37
rect 8811 -62 8857 -47
rect 8737 -5921 8759 -62
rect 8737 -6063 8777 -5921
rect 8817 -5921 8857 -62
rect 21649 -112 21689 -47
rect 21723 -112 21769 -37
rect 14678 -217 14812 -216
rect 8978 -237 14812 -217
rect 8978 -288 9274 -237
rect 14514 -264 14812 -237
rect 14514 -288 14726 -264
rect 8978 -313 14726 -288
rect 8978 -4636 9074 -313
rect 14607 -4634 14726 -313
rect 14542 -4636 14726 -4634
rect 8978 -4680 14726 -4636
rect 14786 -4680 14812 -264
rect 16067 -335 18520 -318
rect 16067 -385 16265 -335
rect 18348 -336 18520 -335
rect 18348 -340 21428 -336
rect 18348 -385 19156 -340
rect 16067 -390 19156 -385
rect 21239 -390 21428 -340
rect 16067 -425 21428 -390
rect 16067 -1724 16174 -425
rect 18413 -442 21428 -425
rect 18413 -1724 18520 -442
rect 16067 -1805 18520 -1724
rect 18961 -443 21428 -442
rect 18961 -1731 19068 -443
rect 21321 -1731 21428 -443
rect 18961 -1805 21428 -1731
rect 16067 -1831 21428 -1805
rect 16070 -1838 21428 -1831
rect 16070 -1844 21427 -1838
rect 16070 -1945 21427 -1935
rect 16070 -1952 21430 -1945
rect 16067 -1978 21430 -1952
rect 16067 -2059 18525 -1978
rect 16067 -4332 16174 -2059
rect 18418 -4332 18525 -2059
rect 16067 -4413 18525 -4332
rect 18964 -2052 21430 -1978
rect 18964 -4329 19071 -2052
rect 21323 -4329 21430 -2052
rect 18964 -4413 21430 -4329
rect 16067 -4436 21430 -4413
rect 16067 -4439 21427 -4436
rect 16070 -4574 21427 -4439
rect 16070 -4633 16364 -4574
rect 18235 -4633 21427 -4574
rect 16070 -4650 21427 -4633
rect 8978 -4730 14812 -4680
rect 14678 -4731 14812 -4730
rect 9076 -4949 13523 -4849
rect 9076 -5735 9176 -4949
rect 13423 -5735 13523 -4949
rect 16046 -4876 19860 -4769
rect 9076 -5825 13523 -5735
rect 9075 -5835 13523 -5825
rect 13959 -5578 14868 -5478
rect 9075 -5836 13521 -5835
rect 9075 -5872 9110 -5836
rect 13477 -5872 13521 -5836
rect 9075 -5905 13521 -5872
rect 13959 -5869 14059 -5578
rect 8811 -6050 8857 -5921
rect 12353 -5991 13874 -5978
rect 12353 -6038 12470 -5991
rect 13775 -6038 13874 -5991
rect 8811 -6063 12074 -6050
rect 8737 -6104 12074 -6063
rect 8737 -6138 8848 -6104
rect 11958 -6138 12074 -6104
rect 8737 -6174 12074 -6138
rect 8737 -6215 8792 -6174
rect 11802 -6184 12074 -6174
rect 11802 -6215 11999 -6184
rect 8737 -6240 11999 -6215
rect 8623 -6879 11541 -6847
rect 8623 -6908 8659 -6879
rect 8589 -6919 8659 -6908
rect 11414 -6919 11541 -6879
rect 8589 -6951 11541 -6919
rect 11437 -6968 11541 -6951
rect 8589 -7111 11075 -7096
rect 8589 -7196 10970 -7111
rect 8589 -7505 8678 -7196
rect 10966 -7373 10970 -7327
rect 11061 -7373 11075 -7111
rect 10975 -7505 11075 -7373
rect 8589 -7605 11075 -7505
rect 11437 -7761 11466 -6968
rect 11507 -7761 11541 -6968
rect 8589 -7976 8678 -7946
rect 8623 -8932 8678 -7976
rect 9607 -8390 9609 -8387
rect 9643 -8390 9661 -8387
rect 9607 -8404 9666 -8390
rect 9607 -8506 9620 -8404
rect 9660 -8506 9666 -8404
rect 9607 -8517 9666 -8506
rect 9982 -8404 10040 -8390
rect 9982 -8506 9994 -8404
rect 10034 -8506 10040 -8404
rect 9982 -8517 10040 -8506
rect 10258 -8404 10316 -8390
rect 10258 -8506 10270 -8404
rect 10310 -8506 10316 -8404
rect 10258 -8517 10316 -8506
rect 10534 -8404 10592 -8390
rect 10534 -8506 10546 -8404
rect 10586 -8506 10592 -8404
rect 10534 -8517 10592 -8506
rect 10809 -8404 10863 -8390
rect 10809 -8506 10817 -8404
rect 10857 -8506 10863 -8404
rect 10809 -8517 10863 -8506
rect 9607 -8519 9661 -8517
rect 9787 -8597 9865 -8586
rect 9417 -8599 9587 -8597
rect 9417 -8639 9431 -8599
rect 9574 -8639 9587 -8599
rect 9417 -8642 9587 -8639
rect 9787 -8649 9799 -8597
rect 9852 -8649 9865 -8597
rect 9787 -8660 9865 -8649
rect 10069 -8597 10141 -8586
rect 10069 -8649 10075 -8597
rect 10128 -8649 10141 -8597
rect 10069 -8660 10141 -8649
rect 10346 -8597 10417 -8586
rect 10346 -8649 10351 -8597
rect 10404 -8649 10417 -8597
rect 10346 -8660 10417 -8649
rect 10622 -8597 10693 -8586
rect 10622 -8649 10627 -8597
rect 10680 -8649 10693 -8597
rect 10622 -8660 10693 -8649
rect 11437 -8880 11462 -7761
rect 11514 -8880 11541 -7761
rect 11437 -8916 11466 -8880
rect 11507 -8916 11541 -8880
rect 11437 -8932 11541 -8916
rect 8623 -8937 11541 -8932
rect 8651 -8960 11541 -8937
rect 8651 -9000 8698 -8960
rect 11453 -9000 11541 -8960
rect 8651 -9036 11541 -9000
rect 8651 -19751 8678 -9036
rect 11952 -9492 11999 -6240
rect 8857 -9493 11999 -9492
rect 8623 -19824 8678 -19751
rect 8737 -9514 11999 -9493
rect 8737 -19631 8761 -9514
rect 8819 -9527 11999 -9514
rect 12033 -9492 12074 -6184
rect 12353 -6078 13874 -6038
rect 12353 -6118 12453 -6078
rect 12353 -8412 12362 -6118
rect 12403 -8345 12453 -6118
rect 13774 -8345 13874 -6078
rect 13959 -7902 13968 -5869
rect 14004 -7840 14059 -5869
rect 14768 -7840 14868 -5578
rect 14004 -7902 14868 -7840
rect 13959 -7940 14868 -7902
rect 12403 -8412 13874 -8345
rect 12353 -8445 13874 -8412
rect 16046 -8743 16153 -4876
rect 18967 -6162 19074 -4876
rect 19753 -4968 19860 -4876
rect 19753 -5075 21266 -4968
rect 19753 -6162 19860 -5075
rect 18967 -6269 19860 -6162
rect 18967 -6316 19268 -6269
rect 18967 -7244 19122 -6316
rect 19215 -7244 19268 -6316
rect 19753 -6609 19860 -6269
rect 18967 -7311 19268 -7244
rect 19614 -6685 19860 -6609
rect 18967 -8743 19074 -7311
rect 16046 -8850 19074 -8743
rect 19614 -8668 19654 -6685
rect 19724 -8668 19860 -6685
rect 21159 -7335 21266 -5075
rect 19614 -8747 19860 -8668
rect 12033 -9527 12077 -9492
rect 8819 -9566 12077 -9527
rect 8819 -9600 8833 -9566
rect 11943 -9600 12077 -9566
rect 8819 -9640 12077 -9600
rect 8819 -19631 8857 -9640
rect 9239 -9898 14177 -9792
rect 9239 -9926 9432 -9898
rect 9239 -9994 9373 -9926
rect 13966 -9926 14177 -9898
rect 9239 -10668 9336 -9994
rect 9370 -10668 9373 -9994
rect 9239 -10738 9373 -10668
rect 14043 -10738 14177 -9926
rect 19753 -9832 19860 -8747
rect 21126 -7433 21266 -7335
rect 21126 -9832 21233 -7433
rect 19753 -9939 21233 -9832
rect 21649 -9259 21679 -112
rect 21731 -9259 21769 -112
rect 9239 -10746 14177 -10738
rect 9239 -10872 14276 -10746
rect 9239 -10960 9373 -10872
rect 14043 -10880 14276 -10872
rect 9239 -11868 9336 -10960
rect 9370 -11868 9373 -10960
rect 9239 -11929 9373 -11868
rect 14142 -11904 14276 -10880
rect 15393 -11044 18497 -11021
rect 15393 -11118 16163 -11044
rect 18451 -11118 18497 -11044
rect 15393 -11193 18497 -11118
rect 15393 -11533 15565 -11193
rect 18325 -11533 18497 -11193
rect 15393 -11583 18497 -11533
rect 14142 -11929 14328 -11904
rect 9239 -12063 14328 -11929
rect 9239 -12120 9373 -12063
rect 9239 -15368 9336 -12120
rect 9370 -15368 9373 -12120
rect 9239 -15461 9373 -15368
rect 14194 -12727 14328 -12063
rect 14194 -15460 14233 -12727
rect 14284 -15460 14328 -12727
rect 15393 -13175 15474 -11583
rect 15532 -11596 18497 -11583
rect 15532 -11647 15644 -11596
rect 18331 -11605 18497 -11596
rect 21649 -11392 21689 -9259
rect 21723 -11392 21769 -9259
rect 18331 -11647 18762 -11605
rect 15532 -11705 18762 -11647
rect 15532 -11772 16874 -11705
rect 15532 -13059 15565 -11772
rect 16702 -13059 16874 -11772
rect 15532 -13175 16874 -13059
rect 15393 -13231 16874 -13175
rect 17297 -11773 18762 -11705
rect 17297 -11777 18664 -11773
rect 17297 -13066 17469 -11777
rect 18590 -13066 18664 -11777
rect 17297 -13198 18664 -13066
rect 18709 -13198 18762 -11773
rect 17297 -13238 18762 -13198
rect 18866 -11701 19670 -11668
rect 18866 -11840 20400 -11701
rect 18866 -12631 19038 -11840
rect 19498 -11873 20400 -11840
rect 19498 -11935 19752 -11873
rect 19498 -12631 19630 -11935
rect 18866 -12858 19630 -12631
rect 14194 -15461 14328 -15460
rect 9239 -15520 14328 -15461
rect 9239 -15578 12233 -15520
rect 14173 -15578 14328 -15520
rect 9239 -15595 14328 -15578
rect 15407 -13375 16905 -13314
rect 11897 -15703 14243 -15647
rect 11897 -15812 14129 -15703
rect 9199 -15885 9364 -15883
rect 9199 -16050 11803 -15885
rect 9199 -17331 9364 -16050
rect 11638 -17331 11803 -16050
rect 9199 -17418 11803 -17331
rect 9199 -17481 10548 -17418
rect 11572 -17481 11803 -17418
rect 9199 -17496 11803 -17481
rect 11897 -17523 12062 -15812
rect 11897 -17529 12070 -17523
rect 14078 -17529 14129 -15812
rect 11897 -17557 14129 -17529
rect 11899 -17586 14129 -17557
rect 11899 -17635 12180 -17586
rect 13979 -17635 14129 -17586
rect 11899 -17694 14129 -17635
rect 9197 -17783 9362 -17781
rect 9197 -17806 11787 -17783
rect 9197 -17869 10546 -17806
rect 11570 -17869 11787 -17806
rect 9197 -17948 11787 -17869
rect 9197 -19225 9362 -17948
rect 11622 -18409 11787 -17948
rect 11622 -19225 11713 -18409
rect 9197 -19356 11713 -19225
rect 11769 -19356 11787 -18409
rect 9197 -19390 11787 -19356
rect 11899 -18418 12070 -17694
rect 11899 -19365 11917 -18418
rect 11973 -19365 12070 -18418
rect 11899 -19406 12070 -19365
rect 14056 -19318 14129 -17694
rect 14191 -17694 14243 -15703
rect 15407 -15828 15479 -13375
rect 15534 -13486 16905 -13375
rect 15534 -15828 15579 -13486
rect 15407 -15852 15579 -15828
rect 16733 -15852 16905 -13486
rect 15407 -16024 16905 -15852
rect 17309 -13482 18810 -13310
rect 17309 -15837 17481 -13482
rect 18638 -13820 18810 -13482
rect 18638 -15821 18705 -13820
rect 18756 -15821 18810 -13820
rect 18866 -14153 19038 -12858
rect 19498 -13572 19630 -12858
rect 19706 -13572 19752 -11935
rect 19498 -13767 19752 -13572
rect 20228 -13767 20400 -11873
rect 19498 -13939 20400 -13767
rect 19498 -14153 19670 -13939
rect 18866 -14325 19670 -14153
rect 18638 -15837 18810 -15821
rect 17309 -16009 18810 -15837
rect 18909 -15003 21549 -14921
rect 18909 -15086 21464 -15003
rect 18909 -15246 19074 -15086
rect 15400 -17171 18833 -17006
rect 14191 -19318 14227 -17694
rect 14056 -19406 14227 -19318
rect 11899 -19577 14227 -19406
rect 15400 -19421 15565 -17171
rect 16875 -19421 17015 -17171
rect 17214 -19421 17354 -17171
rect 18668 -19421 18833 -17171
rect 15400 -19510 18833 -19421
rect 15400 -19567 15772 -19510
rect 18452 -19567 18833 -19510
rect 18909 -19074 18931 -15246
rect 18991 -19074 19074 -15246
rect 18909 -19368 19074 -19074
rect 21384 -19179 21464 -15086
rect 21526 -19179 21549 -15003
rect 21384 -19368 21549 -19179
rect 18909 -19533 21549 -19368
rect 15400 -19586 18833 -19567
rect 8737 -19663 8777 -19631
rect 8811 -19650 8857 -19631
rect 21649 -19612 21677 -11392
rect 21725 -19612 21769 -11392
rect 21649 -19650 21689 -19612
rect 8811 -19663 21689 -19650
rect 21723 -19663 21769 -19612
rect 8737 -19678 21769 -19663
rect 8737 -19689 8877 -19678
rect 21631 -19689 21769 -19678
rect 8737 -19723 8837 -19689
rect 21663 -19723 21769 -19689
rect 8737 -19730 8877 -19723
rect 21631 -19730 21769 -19723
rect 8737 -19755 21769 -19730
rect 21837 -9655 21860 108
rect 21837 -11310 21887 -9655
rect 21837 -19824 21860 -11310
rect 8623 -19837 21860 -19824
rect 8589 -19878 8619 -19843
rect 21812 -19863 21860 -19837
rect 21900 -19863 21921 -19843
rect 21812 -19869 21921 -19863
rect 8589 -19903 8649 -19878
rect 21861 -19903 21921 -19869
<< viali >>
rect 8715 172 21727 178
rect 8715 132 21727 172
rect 8609 -6093 8623 36
rect 8623 -6093 8651 36
rect 8869 23 21623 34
rect 8869 -11 21623 23
rect 8869 -18 21623 -11
rect 8759 -5921 8777 -62
rect 8777 -6063 8811 -62
rect 8811 -5921 8817 -62
rect 9274 -288 14514 -237
rect 14726 -4680 14786 -264
rect 16265 -385 18348 -335
rect 19156 -390 21239 -340
rect 16364 -4633 18235 -4574
rect 9110 -5872 13477 -5836
rect 12470 -6038 13775 -5991
rect 8792 -6215 11802 -6174
rect 10970 -7373 11061 -7111
rect 10033 -7966 10072 -7858
rect 10217 -7966 10256 -7858
rect 10401 -7966 10440 -7858
rect 10585 -7966 10624 -7858
rect 10769 -7966 10808 -7858
rect 9620 -8506 9660 -8404
rect 9994 -8506 10034 -8404
rect 10270 -8506 10310 -8404
rect 10546 -8506 10586 -8404
rect 10817 -8506 10857 -8404
rect 9431 -8639 9574 -8599
rect 9799 -8649 9852 -8597
rect 10075 -8649 10128 -8597
rect 10351 -8649 10404 -8597
rect 10627 -8649 10680 -8597
rect 11462 -8880 11466 -7761
rect 11466 -8880 11507 -7761
rect 11507 -8880 11514 -7761
rect 8609 -19751 8623 -8937
rect 8623 -19751 8651 -8937
rect 8761 -9678 8819 -9514
rect 12362 -8412 12403 -6118
rect 13968 -7902 14004 -5869
rect 19122 -7244 19215 -6316
rect 19654 -8668 19724 -6685
rect 8761 -19631 8777 -9678
rect 8777 -19631 8811 -9678
rect 8811 -19631 8819 -9678
rect 9432 -9932 13966 -9898
rect 9336 -10668 9370 -9994
rect 21679 -9259 21689 -112
rect 21689 -9259 21723 -112
rect 21723 -9259 21731 -112
rect 9336 -11868 9370 -10960
rect 16163 -11118 18451 -11044
rect 9336 -15368 9370 -12120
rect 14233 -15460 14284 -12727
rect 15474 -13175 15532 -11583
rect 15644 -11647 18331 -11596
rect 18664 -13198 18709 -11773
rect 12233 -15578 14173 -15520
rect 10548 -17481 11572 -17418
rect 12180 -17635 13979 -17586
rect 10546 -17869 11570 -17806
rect 11713 -19356 11769 -18409
rect 11917 -19365 11973 -18418
rect 14129 -19318 14191 -15703
rect 15479 -15828 15534 -13375
rect 18705 -15821 18756 -13820
rect 19630 -13572 19706 -11935
rect 15772 -19567 18452 -19510
rect 18931 -19074 18991 -15246
rect 21464 -19179 21526 -15003
rect 21677 -19612 21689 -11392
rect 21689 -19612 21723 -11392
rect 21723 -19612 21725 -11392
rect 8877 -19689 21631 -19678
rect 8877 -19723 21631 -19689
rect 8877 -19730 21631 -19723
rect 21860 -9655 21887 139
rect 21887 -9655 21900 139
rect 8619 -19843 8623 -19837
rect 8623 -19843 21812 -19837
rect 8619 -19869 21812 -19843
rect 21860 -19843 21887 -11310
rect 21887 -19843 21900 -11310
rect 21860 -19863 21900 -19843
rect 8619 -19878 8649 -19869
rect 8649 -19878 21812 -19869
<< metal1 >>
rect 8589 178 21921 206
rect 8589 132 8715 178
rect 21727 139 21921 178
rect 21727 132 21860 139
rect 8589 108 21860 132
rect 8589 36 8678 108
rect 8589 -6093 8609 36
rect 8651 -6093 8678 36
rect 8589 -6122 8678 -6093
rect 8720 34 21780 80
rect 8720 -18 8869 34
rect 21623 -18 21780 34
rect 8720 -62 21780 -18
rect 8720 -5921 8759 -62
rect 8817 -112 21780 -62
rect 8817 -120 21679 -112
rect 8817 -5921 8920 -120
rect 9219 -237 21495 -200
rect 9219 -288 9274 -237
rect 14514 -264 21495 -237
rect 14514 -288 14726 -264
rect 9219 -400 14726 -288
rect 9068 -4238 9132 -450
rect 9219 -2449 11719 -2443
rect 9219 -2501 9225 -2449
rect 11713 -2501 11719 -2449
rect 9219 -2507 11719 -2501
rect 9068 -4482 9074 -4238
rect 9126 -4482 9132 -4238
rect 9068 -4488 9132 -4482
rect 11805 -4250 11869 -450
rect 11955 -2449 14455 -2443
rect 11955 -2501 11961 -2449
rect 14449 -2501 14455 -2449
rect 11955 -2507 14455 -2501
rect 11805 -4494 11811 -4250
rect 11863 -4494 11869 -4250
rect 14542 -4238 14606 -450
rect 14542 -4482 14548 -4238
rect 14600 -4482 14606 -4238
rect 14542 -4488 14606 -4482
rect 11805 -4500 11869 -4494
rect 9219 -4620 11719 -4556
rect 11955 -4620 14455 -4556
rect 14700 -4620 14726 -400
rect 9220 -4680 14726 -4620
rect 14786 -335 21495 -264
rect 14786 -385 16265 -335
rect 18348 -340 21495 -335
rect 18348 -385 19156 -340
rect 14786 -390 19156 -385
rect 21239 -390 21495 -340
rect 14786 -400 21495 -390
rect 14786 -3400 14900 -400
rect 15500 -1700 16000 -1500
rect 15500 -3400 15700 -1700
rect 14786 -3600 15700 -3400
rect 14786 -4680 14900 -3600
rect 15000 -3700 15200 -3694
rect 15200 -3900 15400 -3700
rect 15000 -3906 15400 -3900
rect 15200 -4280 15400 -3906
rect 15180 -4300 15420 -4280
rect 15180 -4500 15200 -4300
rect 15400 -4500 15420 -4300
rect 15180 -4520 15420 -4500
rect 9220 -4820 14900 -4680
rect 14877 -4899 15117 -4878
rect 14877 -4900 14900 -4899
rect 9300 -5012 14900 -4900
rect 8999 -5590 9290 -5089
rect 13348 -5400 13412 -5090
rect 13865 -5116 14106 -5097
rect 13865 -5316 13885 -5116
rect 14085 -5184 14106 -5116
rect 14877 -5099 14900 -5012
rect 15100 -4900 15117 -4899
rect 15200 -4900 15400 -4520
rect 15100 -5099 15400 -4900
rect 14877 -5100 15400 -5099
rect 14877 -5122 15117 -5100
rect 15167 -5175 15428 -5158
rect 15167 -5184 15179 -5175
rect 14085 -5296 15179 -5184
rect 14085 -5316 14106 -5296
rect 13865 -5340 14106 -5316
rect 15167 -5306 15179 -5296
rect 15413 -5306 15428 -5175
rect 15167 -5323 15428 -5306
rect 15180 -5400 15420 -5380
rect 13348 -5590 15200 -5400
rect 8720 -6063 8777 -5921
rect 8811 -6063 8920 -5921
rect 9000 -5800 9200 -5590
rect 13400 -5600 15200 -5590
rect 15400 -5600 15420 -5400
rect 14210 -5652 14610 -5600
rect 15180 -5620 15420 -5600
rect 9300 -5732 14178 -5668
rect 9000 -5836 12100 -5800
rect 12300 -5835 14009 -5800
rect 12300 -5836 14011 -5835
rect 9000 -5872 9110 -5836
rect 13477 -5842 14011 -5836
rect 13477 -5872 13930 -5842
rect 13985 -5869 14011 -5842
rect 9000 -6000 12100 -5872
rect 12300 -5905 13930 -5872
rect 12300 -6000 12306 -5905
rect 12426 -5991 13837 -5975
rect 8720 -6099 8920 -6063
rect 12426 -6038 12470 -5991
rect 13775 -6038 13837 -5991
rect 12426 -6088 13837 -6038
rect 11644 -6099 13837 -6088
rect 8720 -6118 13837 -6099
rect 8720 -6174 12362 -6118
rect 8720 -6215 8792 -6174
rect 11802 -6215 12362 -6174
rect 8720 -6299 12362 -6215
rect 8720 -6300 9065 -6299
rect 11644 -6328 12362 -6299
rect 8589 -6438 8788 -6370
rect 8589 -6446 9057 -6438
rect 8589 -6500 8887 -6446
rect 9041 -6500 9057 -6446
rect 8589 -6506 9057 -6500
rect 8589 -6570 8788 -6506
rect 8589 -6726 8788 -6649
rect 8589 -6734 9056 -6726
rect 8589 -6788 8886 -6734
rect 9040 -6788 9056 -6734
rect 8589 -6794 9056 -6788
rect 8589 -6849 8788 -6794
rect 8706 -6951 10917 -6946
rect 8706 -7012 8714 -6951
rect 8770 -7011 10852 -6951
rect 10908 -7011 10917 -6951
rect 8770 -7012 10917 -7011
rect 8706 -7017 10917 -7012
rect 8591 -7278 10808 -7078
rect 10955 -7111 11075 -7095
rect 8709 -7326 8775 -7319
rect 8709 -7378 8716 -7326
rect 8768 -7378 8775 -7326
rect 8709 -7385 8775 -7378
rect 10847 -7325 10913 -7319
rect 10847 -7377 10854 -7325
rect 10906 -7377 10913 -7325
rect 10847 -7385 10913 -7377
rect 10955 -7373 10970 -7111
rect 11061 -7316 11075 -7111
rect 11191 -7311 11359 -7301
rect 11191 -7316 11203 -7311
rect 11061 -7370 11203 -7316
rect 11348 -7370 11359 -7311
rect 11061 -7373 11359 -7370
rect 10955 -7381 11359 -7373
rect 11644 -7434 11912 -6328
rect 8589 -7705 8789 -7563
rect 8850 -7674 11912 -7434
rect 8589 -7713 9143 -7705
rect 8589 -7763 8973 -7713
rect 8958 -7767 8973 -7763
rect 9127 -7767 9143 -7713
rect 8958 -7773 9143 -7767
rect 10919 -7761 11542 -7721
rect 10919 -7817 11462 -7761
rect 8588 -7887 8788 -7836
rect 10027 -7858 10078 -7845
rect 10027 -7879 10033 -7858
rect 8588 -7900 9144 -7887
rect 8588 -7954 8974 -7900
rect 9128 -7954 9144 -7900
rect 8588 -7964 9144 -7954
rect 9292 -7916 10033 -7879
rect 8588 -8036 8788 -7964
rect 9292 -8112 9329 -7916
rect 10027 -7966 10033 -7916
rect 10072 -7966 10078 -7858
rect 10211 -7858 10262 -7845
rect 10211 -7926 10217 -7858
rect 10027 -7978 10078 -7966
rect 10118 -7964 10217 -7926
rect 8589 -8187 8788 -8121
rect 8980 -8149 9329 -8112
rect 9609 -8036 9677 -8021
rect 8980 -8187 9017 -8149
rect 8589 -8200 9017 -8187
rect 8589 -8254 8830 -8200
rect 8984 -8254 9017 -8200
rect 9609 -8190 9615 -8036
rect 9669 -8190 9677 -8036
rect 9609 -8206 9677 -8190
rect 9812 -8031 9880 -8020
rect 10118 -8031 10156 -7964
rect 10211 -7966 10217 -7964
rect 10256 -7966 10262 -7858
rect 10395 -7858 10446 -7845
rect 10395 -7924 10401 -7858
rect 10211 -7978 10262 -7966
rect 10290 -7964 10401 -7924
rect 9812 -8035 10156 -8031
rect 9812 -8189 9818 -8035
rect 9872 -8069 10156 -8035
rect 10185 -8030 10253 -8018
rect 10290 -8030 10330 -7964
rect 10395 -7966 10401 -7964
rect 10440 -7966 10446 -7858
rect 10579 -7858 10630 -7845
rect 10579 -7897 10585 -7858
rect 10395 -7978 10446 -7966
rect 10543 -7966 10585 -7897
rect 10624 -7966 10630 -7858
rect 10543 -7978 10630 -7966
rect 10763 -7858 10814 -7845
rect 10763 -7966 10769 -7858
rect 10808 -7966 10814 -7858
rect 10763 -7978 10814 -7966
rect 10185 -8033 10330 -8030
rect 9872 -8189 9880 -8069
rect 9812 -8205 9880 -8189
rect 10185 -8187 10191 -8033
rect 10245 -8070 10330 -8033
rect 10365 -8028 10433 -8013
rect 10245 -8187 10253 -8070
rect 10185 -8203 10253 -8187
rect 10365 -8182 10371 -8028
rect 10425 -8030 10433 -8028
rect 10543 -8030 10583 -7978
rect 10425 -8070 10583 -8030
rect 10636 -8028 10704 -8013
rect 10425 -8182 10433 -8070
rect 10365 -8198 10433 -8182
rect 10636 -8182 10642 -8028
rect 10696 -8029 10704 -8028
rect 10765 -8029 10805 -7978
rect 10696 -8069 10805 -8029
rect 10696 -8182 10704 -8069
rect 10636 -8198 10704 -8182
rect 8589 -8264 9017 -8254
rect 8589 -8321 8788 -8264
rect 11108 -8265 11344 -8261
rect 9126 -8361 9411 -8265
rect 10963 -8269 11344 -8265
rect 10963 -8354 11118 -8269
rect 11331 -8354 11344 -8269
rect 10963 -8361 11344 -8354
rect 8590 -8453 8790 -8400
rect 9126 -8453 9222 -8361
rect 11108 -8363 11344 -8361
rect 8590 -8549 9222 -8453
rect 9608 -8393 9672 -8390
rect 9608 -8511 9614 -8393
rect 9666 -8511 9672 -8393
rect 9608 -8517 9672 -8511
rect 9982 -8404 10040 -8390
rect 9982 -8459 9994 -8404
rect 10034 -8453 10040 -8404
rect 10258 -8404 10316 -8390
rect 10258 -8452 10270 -8404
rect 10034 -8459 10046 -8453
rect 9982 -8511 9988 -8459
rect 10040 -8511 10046 -8459
rect 9982 -8517 10046 -8511
rect 10257 -8458 10270 -8452
rect 10310 -8452 10316 -8404
rect 10534 -8404 10592 -8390
rect 10310 -8458 10321 -8452
rect 10534 -8453 10546 -8404
rect 10257 -8510 10263 -8458
rect 10315 -8510 10321 -8458
rect 10257 -8516 10321 -8510
rect 10533 -8458 10546 -8453
rect 10586 -8453 10592 -8404
rect 10805 -8404 10863 -8390
rect 10586 -8458 10597 -8453
rect 10533 -8511 10539 -8458
rect 10591 -8511 10597 -8458
rect 10258 -8518 10316 -8516
rect 10533 -8517 10597 -8511
rect 10805 -8458 10817 -8404
rect 10857 -8453 10863 -8404
rect 10857 -8458 10869 -8453
rect 10805 -8511 10810 -8458
rect 10863 -8511 10869 -8458
rect 10805 -8517 10869 -8511
rect 10534 -8518 10592 -8517
rect 8590 -8600 8790 -8549
rect 9411 -8592 9596 -8584
rect 9411 -8646 9426 -8592
rect 9574 -8603 9596 -8592
rect 9787 -8597 9865 -8586
rect 9574 -8640 9597 -8603
rect 9574 -8646 9596 -8640
rect 9411 -8652 9596 -8646
rect 9787 -8649 9799 -8597
rect 9852 -8649 9865 -8597
rect 9787 -8660 9865 -8649
rect 10063 -8597 10141 -8586
rect 10063 -8649 10075 -8597
rect 10128 -8649 10141 -8597
rect 10063 -8660 10141 -8649
rect 10339 -8597 10417 -8586
rect 10339 -8649 10351 -8597
rect 10404 -8649 10417 -8597
rect 10339 -8660 10417 -8649
rect 10615 -8597 10693 -8586
rect 10615 -8649 10627 -8597
rect 10680 -8649 10693 -8597
rect 10615 -8660 10693 -8649
rect 8587 -8809 8790 -8705
rect 11434 -8809 11462 -7817
rect 8587 -8880 11462 -8809
rect 11514 -8880 11542 -7761
rect 8587 -8905 11542 -8880
rect 11644 -8600 11912 -7674
rect 12283 -8412 12362 -6328
rect 12403 -6158 13837 -6118
rect 12403 -8412 12412 -6158
rect 12468 -6214 12532 -6208
rect 12468 -8194 12474 -6214
rect 12526 -8194 12532 -6214
rect 12468 -8200 12532 -8194
rect 13706 -6214 13770 -6208
rect 13706 -8194 13712 -6214
rect 13764 -8194 13770 -6214
rect 13903 -7958 13930 -5905
rect 14004 -7902 14011 -5869
rect 13985 -7958 14011 -7902
rect 13903 -8001 14011 -7958
rect 14068 -7756 14132 -5732
rect 14688 -7756 14752 -5708
rect 15500 -6611 15700 -3600
rect 15800 -4000 16000 -1800
rect 15800 -4206 16000 -4200
rect 15800 -4300 16000 -4294
rect 15800 -4506 16000 -4500
rect 15786 -4574 18257 -4562
rect 15786 -4633 16364 -4574
rect 18235 -4633 18257 -4574
rect 15786 -4681 18257 -4633
rect 15786 -5156 15985 -4681
rect 15760 -5170 16018 -5156
rect 15760 -5301 15772 -5170
rect 16006 -5301 16018 -5170
rect 15760 -5316 16018 -5301
rect 15780 -5400 16020 -5380
rect 15780 -5600 15800 -5400
rect 16000 -5600 16020 -5400
rect 15780 -5620 16020 -5600
rect 15499 -6803 15700 -6611
rect 14068 -7800 14752 -7756
rect 14068 -8000 14900 -7800
rect 15100 -8000 15106 -7800
rect 13706 -8200 13770 -8194
rect 12619 -8300 13619 -8256
rect 15180 -8300 15420 -8280
rect 12619 -8352 15200 -8300
rect 12283 -8439 12412 -8412
rect 12700 -8500 15200 -8352
rect 15400 -8500 15420 -8300
rect 15180 -8520 15420 -8500
rect 14580 -8600 14820 -8580
rect 15500 -8600 15700 -6803
rect 11644 -8800 14600 -8600
rect 14800 -8800 15700 -8600
rect 11644 -8897 15700 -8800
rect 15800 -8700 16000 -5620
rect 19074 -6316 19270 -6261
rect 19074 -7244 19122 -6316
rect 19215 -7118 19270 -6316
rect 19614 -6685 19757 -6609
rect 19614 -7118 19654 -6685
rect 19215 -7244 19654 -7118
rect 19074 -7314 19654 -7244
rect 19614 -8668 19654 -7314
rect 19724 -8668 19757 -6685
rect 19614 -8679 19757 -8668
rect 8588 -8937 8677 -8905
rect 8588 -9040 8609 -8937
rect 8589 -19751 8609 -9040
rect 8651 -9018 8677 -8937
rect 11644 -9017 11912 -8897
rect 15800 -8900 19000 -8700
rect 19200 -8900 19206 -8700
rect 8651 -19751 8678 -9018
rect 8589 -19824 8678 -19751
rect 8720 -9223 11912 -9017
rect 8720 -9514 8920 -9223
rect 10234 -9296 10298 -9290
rect 10234 -9330 10240 -9296
rect 8720 -19631 8761 -9514
rect 8819 -19580 8920 -9514
rect 9060 -9348 10240 -9330
rect 10292 -9348 10298 -9296
rect 9060 -9354 10298 -9348
rect 9060 -9390 10296 -9354
rect 9060 -17772 9120 -9390
rect 10820 -9450 10880 -9444
rect 9180 -9510 10820 -9450
rect 14280 -9500 14520 -9480
rect 19600 -9482 19800 -8679
rect 21580 -9101 21679 -120
rect 21314 -9301 21320 -9101
rect 21520 -9259 21679 -9101
rect 21731 -9259 21780 -112
rect 21520 -9301 21780 -9259
rect 19578 -9500 19811 -9482
rect 9180 -15770 9240 -9510
rect 10820 -9516 10880 -9510
rect 12080 -9595 12100 -9500
rect 9300 -9700 12100 -9595
rect 12300 -9700 14300 -9500
rect 14500 -9700 19600 -9500
rect 19800 -9700 19811 -9500
rect 21837 -9655 21860 108
rect 21900 -9655 21921 139
rect 21837 -9700 21921 -9655
rect 9300 -9880 14100 -9700
rect 14280 -9720 14520 -9700
rect 19578 -9721 19811 -9700
rect 9300 -9898 14098 -9880
rect 9300 -9932 9432 -9898
rect 13966 -9932 14098 -9898
rect 9300 -9938 14098 -9932
rect 9300 -9994 9376 -9938
rect 9300 -10668 9336 -9994
rect 9370 -10668 9376 -9994
rect 15194 -10000 15200 -9800
rect 15400 -10000 18700 -9800
rect 18900 -10000 18906 -9800
rect 18994 -10000 19000 -9800
rect 19200 -9867 19805 -9800
rect 21357 -9867 21910 -9800
rect 19200 -10000 21910 -9867
rect 9471 -10158 13299 -10040
rect 13925 -10100 14300 -10040
rect 13925 -10158 20500 -10100
rect 13199 -10274 13299 -10158
rect 9471 -10626 9892 -10274
rect 13199 -10392 13925 -10274
rect 14100 -10300 20500 -10158
rect 20700 -10300 21910 -10100
rect 17880 -10400 18120 -10380
rect 14100 -10508 17900 -10400
rect 13925 -10600 17900 -10508
rect 18100 -10600 21910 -10400
rect 13925 -10626 14300 -10600
rect 17880 -10620 18120 -10600
rect 9300 -10960 9376 -10668
rect 9300 -11868 9336 -10960
rect 9370 -11868 9376 -10960
rect 14100 -10900 21910 -10700
rect 14100 -11004 14220 -10900
rect 9472 -11356 9893 -11004
rect 13597 -11122 14220 -11004
rect 9472 -11824 9893 -11472
rect 13592 -11600 14024 -11228
rect 15458 -11558 15596 -11021
rect 15800 -11400 16000 -10900
rect 18396 -11010 21910 -11000
rect 16127 -11044 21910 -11010
rect 16127 -11118 16163 -11044
rect 18451 -11076 21910 -11044
rect 18451 -11118 19600 -11076
rect 16127 -11133 19600 -11118
rect 18393 -11200 19600 -11133
rect 17894 -11500 17900 -11300
rect 18100 -11500 18106 -11300
rect 18393 -11558 18551 -11200
rect 15458 -11583 18551 -11558
rect 14018 -11824 14220 -11706
rect 9300 -12120 9376 -11868
rect 9300 -15368 9336 -12120
rect 9370 -15368 9376 -12120
rect 14100 -12164 14220 -11824
rect 9472 -12516 9893 -12164
rect 13651 -12282 14000 -12164
rect 14072 -12282 15400 -12164
rect 9472 -12984 9893 -12632
rect 13651 -12750 14072 -12398
rect 14211 -12727 14300 -12700
rect 9472 -13452 9893 -13100
rect 13651 -13218 14072 -12866
rect 9472 -13920 9893 -13568
rect 13651 -13686 14072 -13334
rect 9472 -14388 9893 -14036
rect 13651 -14154 14072 -13802
rect 9472 -14856 9893 -14504
rect 13651 -14622 14072 -14270
rect 9472 -15324 9893 -14972
rect 13651 -15090 14072 -14738
rect 11700 -15324 13772 -15206
rect 9300 -15500 9376 -15368
rect 11700 -15700 11900 -15324
rect 14211 -15460 14233 -12727
rect 14284 -12900 14300 -12727
rect 14500 -12900 14506 -12700
rect 14594 -12900 14600 -12700
rect 14800 -12900 14806 -12700
rect 14894 -12900 14900 -12700
rect 15100 -12900 15106 -12700
rect 14284 -15460 14500 -12900
rect 14211 -15500 14500 -15460
rect 12200 -15520 14500 -15500
rect 12200 -15578 12233 -15520
rect 14173 -15578 14500 -15520
rect 12200 -15700 14500 -15578
rect 14113 -15703 14500 -15700
rect 9180 -15830 9310 -15770
rect 9280 -17400 9520 -17380
rect 9280 -17600 9300 -17400
rect 9500 -17600 9520 -17400
rect 10547 -17406 10599 -16193
rect 11532 -17406 11584 -16186
rect 9280 -17620 9520 -17600
rect 10527 -17418 11609 -17406
rect 10527 -17481 10548 -17418
rect 11572 -17481 11609 -17418
rect 10527 -17593 11609 -17481
rect 14113 -17568 14129 -15703
rect 12146 -17586 14129 -17568
rect 9060 -17832 9300 -17772
rect 10527 -17806 11606 -17593
rect 12146 -17635 12180 -17586
rect 13979 -17635 14129 -17586
rect 12146 -17664 14129 -17635
rect 10527 -17869 10546 -17806
rect 11570 -17869 11606 -17806
rect 10527 -17884 11606 -17869
rect 11700 -18409 11991 -18379
rect 9280 -19300 9520 -19280
rect 9280 -19500 9300 -19300
rect 9500 -19500 9520 -19300
rect 9280 -19520 9520 -19500
rect 11700 -19356 11713 -18409
rect 11769 -18418 11991 -18409
rect 11769 -19356 11917 -18418
rect 11700 -19365 11917 -19356
rect 11973 -19365 11991 -18418
rect 11700 -19387 11991 -19365
rect 14113 -19318 14129 -17664
rect 14191 -19318 14500 -15703
rect 14600 -16608 14800 -12900
rect 14900 -16308 15100 -12900
rect 15200 -16008 15400 -12282
rect 15458 -13175 15474 -11583
rect 15532 -11596 18551 -11583
rect 15532 -11647 15644 -11596
rect 18331 -11647 18551 -11596
rect 18700 -11350 19300 -11250
rect 18700 -11500 18800 -11350
rect 19200 -11500 19300 -11350
rect 18700 -11600 19300 -11500
rect 19500 -11500 19600 -11200
rect 19800 -11200 21910 -11076
rect 19800 -11500 19900 -11200
rect 19500 -11600 19900 -11500
rect 20400 -11360 20800 -11260
rect 21837 -11310 21921 -11267
rect 20400 -11560 20500 -11360
rect 20700 -11560 20800 -11360
rect 21314 -11550 21320 -11350
rect 21520 -11392 21780 -11350
rect 21520 -11550 21677 -11392
rect 15532 -11657 18551 -11647
rect 15532 -11674 18727 -11657
rect 15532 -13175 15596 -11674
rect 18394 -11733 18727 -11674
rect 15458 -13375 15596 -13175
rect 15458 -15828 15479 -13375
rect 15534 -15828 15596 -13375
rect 15458 -15865 15596 -15828
rect 18633 -11773 18727 -11733
rect 18633 -13198 18664 -11773
rect 18709 -12681 18727 -11773
rect 18800 -11908 19000 -11600
rect 19600 -11908 19800 -11600
rect 20400 -11660 20800 -11560
rect 20500 -11908 20700 -11660
rect 19610 -11935 19726 -11908
rect 18709 -13198 18765 -12681
rect 18633 -13234 18765 -13198
rect 18633 -13755 18727 -13234
rect 19610 -13572 19630 -11935
rect 19706 -13572 19726 -11935
rect 19610 -13604 19726 -13572
rect 18633 -13820 18785 -13755
rect 18633 -15821 18705 -13820
rect 18756 -15821 18785 -13820
rect 21580 -14706 21677 -11550
rect 18633 -15904 18785 -15821
rect 18913 -15246 19025 -14937
rect 15200 -16208 15700 -16008
rect 14900 -16508 15700 -16308
rect 14600 -16808 15700 -16608
rect 18913 -19074 18931 -15246
rect 18991 -19074 19025 -15246
rect 18913 -19119 19025 -19074
rect 21427 -15003 21677 -14706
rect 21427 -19179 21464 -15003
rect 21526 -19179 21677 -15003
rect 21427 -19229 21677 -19179
rect 14113 -19387 14500 -19318
rect 11700 -19525 14500 -19387
rect 15718 -19510 18520 -19473
rect 15718 -19567 15772 -19510
rect 18452 -19567 18520 -19510
rect 15718 -19580 18520 -19567
rect 21580 -19580 21677 -19229
rect 8819 -19612 21677 -19580
rect 21725 -19612 21780 -11392
rect 8819 -19631 21780 -19612
rect 8720 -19678 21780 -19631
rect 8720 -19730 8877 -19678
rect 21631 -19730 21780 -19678
rect 8720 -19780 21780 -19730
rect 21837 -19824 21860 -11310
rect 8589 -19837 21860 -19824
rect 8589 -19878 8619 -19837
rect 21812 -19863 21860 -19837
rect 21900 -19863 21921 -11310
rect 21812 -19878 21921 -19863
rect 8589 -19903 21921 -19878
<< via1 >>
rect 9225 -2501 11713 -2449
rect 9074 -4482 9126 -4238
rect 11961 -2501 14449 -2449
rect 11811 -4494 11863 -4250
rect 14548 -4482 14600 -4238
rect 15000 -3900 15200 -3700
rect 15200 -4500 15400 -4300
rect 13885 -5316 14085 -5116
rect 14900 -5099 15100 -4899
rect 15179 -5306 15413 -5175
rect 15200 -5600 15400 -5400
rect 12100 -5836 12300 -5800
rect 12100 -5872 12300 -5836
rect 13930 -5869 13985 -5842
rect 12100 -6000 12300 -5872
rect 8887 -6500 9041 -6446
rect 8886 -6788 9040 -6734
rect 8714 -7012 8770 -6951
rect 10852 -7011 10908 -6951
rect 8716 -7378 8768 -7326
rect 10854 -7377 10906 -7325
rect 11203 -7370 11348 -7311
rect 8973 -7767 9127 -7713
rect 8974 -7954 9128 -7900
rect 8830 -8254 8984 -8200
rect 9615 -8190 9669 -8036
rect 9818 -8189 9872 -8035
rect 10191 -8187 10245 -8033
rect 10371 -8182 10425 -8028
rect 10642 -8182 10696 -8028
rect 11118 -8354 11331 -8269
rect 9614 -8404 9666 -8393
rect 9614 -8506 9620 -8404
rect 9620 -8506 9660 -8404
rect 9660 -8506 9666 -8404
rect 9614 -8511 9666 -8506
rect 9988 -8506 9994 -8459
rect 9994 -8506 10034 -8459
rect 10034 -8506 10040 -8459
rect 9988 -8511 10040 -8506
rect 10263 -8506 10270 -8458
rect 10270 -8506 10310 -8458
rect 10310 -8506 10315 -8458
rect 10263 -8510 10315 -8506
rect 10539 -8506 10546 -8458
rect 10546 -8506 10586 -8458
rect 10586 -8506 10591 -8458
rect 10539 -8511 10591 -8506
rect 10810 -8506 10817 -8458
rect 10817 -8506 10857 -8458
rect 10857 -8506 10863 -8458
rect 10810 -8511 10863 -8506
rect 9426 -8599 9574 -8592
rect 9426 -8639 9431 -8599
rect 9431 -8639 9574 -8599
rect 9426 -8646 9574 -8639
rect 9799 -8649 9852 -8597
rect 10075 -8649 10128 -8597
rect 10351 -8649 10404 -8597
rect 10627 -8649 10680 -8597
rect 12474 -8194 12526 -6214
rect 13712 -8194 13764 -6214
rect 13930 -7902 13968 -5869
rect 13968 -7902 13985 -5869
rect 13930 -7958 13985 -7902
rect 15800 -4200 16000 -4000
rect 15800 -4500 16000 -4300
rect 15772 -5301 16006 -5170
rect 15800 -5600 16000 -5400
rect 14900 -8000 15100 -7800
rect 15200 -8500 15400 -8300
rect 14600 -8800 14800 -8600
rect 19000 -8900 19200 -8700
rect 10240 -9348 10292 -9296
rect 10820 -9510 10880 -9450
rect 21320 -9301 21520 -9101
rect 12100 -9700 12300 -9500
rect 14300 -9700 14500 -9500
rect 19600 -9700 19800 -9500
rect 15200 -10000 15400 -9800
rect 18700 -10000 18900 -9800
rect 19000 -10000 19200 -9800
rect 20500 -10300 20700 -10100
rect 17900 -10600 18100 -10400
rect 17900 -11500 18100 -11300
rect 14300 -12900 14500 -12700
rect 14600 -12900 14800 -12700
rect 14900 -12900 15100 -12700
rect 9300 -17600 9500 -17400
rect 9300 -19500 9500 -19300
rect 18800 -11500 19200 -11350
rect 19600 -11500 19800 -11076
rect 20500 -11560 20700 -11360
rect 21320 -11550 21520 -11350
<< metal2 >>
rect 9219 -2449 15200 -2411
rect 9219 -2501 9225 -2449
rect 11713 -2501 11961 -2449
rect 14449 -2501 15200 -2449
rect 9219 -2539 15200 -2501
rect 15000 -3700 15200 -2539
rect 14994 -3900 15000 -3700
rect 15200 -3900 15206 -3700
rect 14900 -4200 15800 -4000
rect 16000 -4200 16006 -4000
rect 9068 -4238 9132 -4232
rect 9068 -4482 9074 -4238
rect 9126 -4482 9132 -4238
rect 14542 -4238 14606 -4232
rect 9068 -4556 9132 -4482
rect 11805 -4250 11869 -4244
rect 11805 -4494 11811 -4250
rect 11863 -4494 11869 -4250
rect 11805 -4556 11869 -4494
rect 14542 -4482 14548 -4238
rect 14600 -4482 14606 -4238
rect 14542 -4556 14606 -4482
rect 14900 -4556 15100 -4200
rect 15180 -4300 15420 -4280
rect 15180 -4500 15200 -4300
rect 15400 -4500 15800 -4300
rect 16000 -4500 16006 -4300
rect 15180 -4520 15420 -4500
rect 9068 -4620 15100 -4556
rect 12100 -5800 12300 -5794
rect 13600 -5800 13770 -4620
rect 14877 -4899 15117 -4878
rect 13865 -5116 14106 -5097
rect 13865 -5316 13885 -5116
rect 14085 -5316 14106 -5116
rect 14877 -5099 14900 -4899
rect 15100 -5099 15117 -4899
rect 14877 -5122 15117 -5099
rect 13865 -5340 14106 -5316
rect 8872 -6445 9057 -6438
rect 8872 -6446 9381 -6445
rect 8872 -6500 8887 -6446
rect 9041 -6493 9381 -6446
rect 9041 -6500 9057 -6493
rect 8872 -6506 9057 -6500
rect 8871 -6734 9056 -6726
rect 8871 -6788 8886 -6734
rect 9040 -6782 9265 -6734
rect 9040 -6788 9056 -6782
rect 8871 -6794 9056 -6788
rect 8709 -6951 8775 -6942
rect 8709 -7012 8714 -6951
rect 8770 -7012 8775 -6951
rect 8709 -7326 8775 -7012
rect 8709 -7378 8716 -7326
rect 8768 -7378 8775 -7326
rect 8709 -7583 8775 -7378
rect 8709 -7662 8913 -7583
rect 8830 -8027 8913 -7662
rect 8958 -7713 9155 -7705
rect 8958 -7767 8973 -7713
rect 9127 -7767 9155 -7713
rect 9217 -7714 9265 -6782
rect 9333 -7607 9381 -6493
rect 10847 -6951 10913 -6943
rect 10847 -7011 10852 -6951
rect 10908 -7011 10913 -6951
rect 10847 -7325 10913 -7011
rect 10847 -7377 10854 -7325
rect 10906 -7377 10913 -7325
rect 9333 -7655 10697 -7607
rect 10847 -7622 10913 -7377
rect 11191 -7311 11359 -7301
rect 11191 -7370 11203 -7311
rect 11348 -7370 11359 -7311
rect 11191 -7381 11359 -7370
rect 9217 -7762 10426 -7714
rect 8958 -7773 9155 -7767
rect 9107 -7810 9155 -7773
rect 9107 -7858 10243 -7810
rect 8959 -7900 9144 -7892
rect 8959 -7954 8974 -7900
rect 9128 -7906 9144 -7900
rect 9128 -7954 9875 -7906
rect 8959 -7960 9144 -7954
rect 9827 -8020 9875 -7954
rect 10195 -8018 10243 -7858
rect 10378 -8013 10426 -7762
rect 10649 -8013 10697 -7655
rect 9609 -8027 9677 -8021
rect 8830 -8036 9677 -8027
rect 8830 -8110 9615 -8036
rect 9609 -8190 9615 -8110
rect 9669 -8190 9677 -8036
rect 8815 -8200 9217 -8192
rect 8815 -8254 8830 -8200
rect 8984 -8254 9217 -8200
rect 9609 -8206 9677 -8190
rect 9812 -8035 9880 -8020
rect 9812 -8189 9818 -8035
rect 9872 -8189 9880 -8035
rect 10185 -8033 10253 -8018
rect 10185 -8152 10191 -8033
rect 9812 -8205 9880 -8189
rect 10097 -8187 10191 -8152
rect 10245 -8187 10253 -8033
rect 8815 -8260 9217 -8254
rect 9149 -8585 9217 -8260
rect 9612 -8387 9672 -8206
rect 9608 -8393 9676 -8387
rect 9608 -8511 9614 -8393
rect 9666 -8511 9676 -8393
rect 9608 -8519 9676 -8511
rect 9411 -8585 9596 -8584
rect 9149 -8592 9598 -8585
rect 9821 -8586 9868 -8205
rect 10097 -8208 10253 -8187
rect 10365 -8028 10433 -8013
rect 10365 -8182 10371 -8028
rect 10425 -8182 10433 -8028
rect 10365 -8198 10433 -8182
rect 10636 -8028 10704 -8013
rect 10636 -8182 10642 -8028
rect 10696 -8182 10704 -8028
rect 10636 -8198 10704 -8182
rect 9149 -8646 9426 -8592
rect 9574 -8646 9598 -8592
rect 9149 -8653 9598 -8646
rect 9787 -8597 9868 -8586
rect 9787 -8649 9799 -8597
rect 9852 -8649 9868 -8597
rect 9787 -8659 9868 -8649
rect 9955 -8459 10051 -8453
rect 9955 -8511 9988 -8459
rect 10040 -8511 10051 -8459
rect 9955 -8514 10051 -8511
rect 9787 -8660 9865 -8659
rect 9955 -9270 10020 -8514
rect 10097 -8586 10144 -8208
rect 10063 -8597 10144 -8586
rect 10063 -8649 10075 -8597
rect 10128 -8649 10144 -8597
rect 10063 -8659 10144 -8649
rect 10231 -8458 10330 -8451
rect 10231 -8510 10263 -8458
rect 10315 -8510 10330 -8458
rect 10231 -8512 10330 -8510
rect 10063 -8660 10141 -8659
rect 9000 -9330 10020 -9270
rect 10231 -9290 10300 -8512
rect 10373 -8586 10420 -8198
rect 10339 -8597 10420 -8586
rect 10339 -8649 10351 -8597
rect 10404 -8649 10420 -8597
rect 10339 -8659 10420 -8649
rect 10507 -8458 10606 -8453
rect 10507 -8511 10539 -8458
rect 10591 -8511 10606 -8458
rect 10507 -8514 10606 -8511
rect 10339 -8660 10417 -8659
rect 10231 -9292 10298 -9290
rect 10234 -9296 10298 -9292
rect 9000 -19369 9060 -9330
rect 10234 -9348 10240 -9296
rect 10292 -9348 10298 -9296
rect 10234 -9354 10298 -9348
rect 10507 -9390 10571 -8514
rect 10649 -8586 10696 -8198
rect 11206 -8261 11343 -7381
rect 11108 -8269 11344 -8261
rect 11108 -8354 11118 -8269
rect 11331 -8354 11344 -8269
rect 11108 -8363 11344 -8354
rect 10805 -8458 10877 -8452
rect 10805 -8511 10810 -8458
rect 10863 -8511 10877 -8458
rect 10805 -8521 10877 -8511
rect 10615 -8597 10696 -8586
rect 10615 -8649 10627 -8597
rect 10680 -8649 10696 -8597
rect 10615 -8659 10696 -8649
rect 10615 -8660 10693 -8659
rect 10813 -9268 10877 -8521
rect 10813 -9389 10880 -9268
rect 9120 -9450 10571 -9390
rect 10820 -9450 10880 -9389
rect 9120 -17470 9180 -9450
rect 10814 -9510 10820 -9450
rect 10880 -9510 10886 -9450
rect 12100 -9500 12300 -6000
rect 12468 -6000 13770 -5800
rect 12468 -6214 12532 -6000
rect 12468 -8194 12474 -6214
rect 12526 -8194 12532 -6214
rect 12468 -8200 12532 -8194
rect 13706 -6214 13770 -6000
rect 13706 -8194 13712 -6214
rect 13764 -8194 13770 -6214
rect 13915 -5842 14034 -5340
rect 13915 -7958 13930 -5842
rect 13985 -7958 14034 -5842
rect 13915 -7982 14034 -7958
rect 14900 -7800 15100 -5122
rect 15167 -5175 15428 -5158
rect 15760 -5170 16018 -5156
rect 15760 -5175 15772 -5170
rect 15167 -5306 15179 -5175
rect 15413 -5301 15772 -5175
rect 16006 -5301 16018 -5170
rect 15413 -5304 16018 -5301
rect 15413 -5306 15428 -5304
rect 15167 -5323 15428 -5306
rect 15760 -5316 16018 -5304
rect 15180 -5400 15420 -5380
rect 15780 -5400 16020 -5380
rect 15180 -5600 15200 -5400
rect 15400 -5600 15800 -5400
rect 16000 -5600 16020 -5400
rect 15180 -5620 15420 -5600
rect 15780 -5620 16020 -5600
rect 13706 -8200 13770 -8194
rect 14580 -8600 14820 -8580
rect 14580 -8800 14600 -8600
rect 14800 -8800 14820 -8600
rect 14580 -8820 14820 -8800
rect 12100 -9706 12300 -9700
rect 14280 -9500 14520 -9480
rect 14280 -9700 14300 -9500
rect 14500 -9700 14520 -9500
rect 14280 -9720 14520 -9700
rect 14300 -12700 14500 -9720
rect 14300 -12906 14500 -12900
rect 14600 -12700 14800 -8820
rect 14600 -12906 14800 -12900
rect 14900 -12700 15100 -8000
rect 15180 -8300 15420 -8280
rect 15180 -8500 15200 -8300
rect 15400 -8500 15420 -8300
rect 15180 -8520 15420 -8500
rect 15200 -9800 15400 -8520
rect 19000 -8700 19200 -8694
rect 15200 -10006 15400 -10000
rect 18700 -9800 18900 -9794
rect 17880 -10400 18120 -10380
rect 17880 -10600 17900 -10400
rect 18100 -10600 18120 -10400
rect 17880 -10620 18120 -10600
rect 17900 -11300 18100 -10620
rect 17900 -11506 18100 -11500
rect 18700 -11250 18900 -10000
rect 19000 -9800 19200 -8900
rect 21320 -9101 21520 -9095
rect 19578 -9500 19816 -9482
rect 19578 -9700 19600 -9500
rect 19800 -9700 19816 -9500
rect 19578 -9721 19816 -9700
rect 19000 -10006 19200 -10000
rect 19600 -11000 19800 -9721
rect 20500 -10100 20700 -10094
rect 19500 -11076 19900 -11000
rect 18700 -11350 19300 -11250
rect 18700 -11500 18800 -11350
rect 19200 -11500 19300 -11350
rect 18700 -11600 19300 -11500
rect 19500 -11500 19600 -11076
rect 19800 -11500 19900 -11076
rect 20500 -11260 20700 -10300
rect 19500 -11600 19900 -11500
rect 20400 -11360 20800 -11260
rect 20400 -11560 20500 -11360
rect 20700 -11560 20800 -11360
rect 21320 -11350 21520 -9301
rect 21320 -11556 21520 -11550
rect 20400 -11660 20800 -11560
rect 14900 -12906 15100 -12900
rect 9280 -17400 9520 -17380
rect 9280 -17470 9300 -17400
rect 9120 -17530 9300 -17470
rect 9280 -17600 9300 -17530
rect 9500 -17600 9520 -17400
rect 9280 -17620 9520 -17600
rect 9280 -19300 9520 -19280
rect 9280 -19369 9300 -19300
rect 9000 -19429 9300 -19369
rect 9280 -19500 9300 -19429
rect 9500 -19500 9520 -19300
rect 9280 -19520 9520 -19500
use sky130_fd_pr__res_xhigh_po_0p69_E9MCU4  R1
timestamp 1713140876
transform 0 1 11699 -1 0 -10331
box -469 -2399 469 2399
use sky130_fd_pr__res_xhigh_po_0p69_39QBTQ  R2
timestamp 1713056482
transform 0 1 16942 -1 0 -11365
box -235 -1442 235 1442
use sky130_fd_pr__res_xhigh_po_0p69_NB3ZKH  R3
timestamp 1713140876
transform 0 1 11745 -1 0 -11414
box -586 -2445 586 2445
use sky130_fd_pr__res_xhigh_po_0p69_GAZAU4  R4
timestamp 1713140876
transform 0 -1 11772 1 0 -13744
box -1756 -2472 1756 2472
use sky130_fd_sc_hd__buf_1  sky130_fd_sc_hd__buf_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1715205430
transform 1 0 10604 0 1 -8857
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  sky130_fd_sc_hd__buf_1_2
timestamp 1715205430
transform 1 0 9776 0 1 -8857
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  sky130_fd_sc_hd__buf_1_3
timestamp 1715205430
transform 1 0 10052 0 1 -8857
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  sky130_fd_sc_hd__buf_1_4
timestamp 1715205430
transform 1 0 10328 0 1 -8857
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1715205430
transform 1 0 9408 0 -1 -7769
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  sky130_fd_sc_hd__diode_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1715205430
transform 1 0 10328 0 -1 -7769
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  sky130_fd_sc_hd__diode_2_1
timestamp 1715205430
transform 1 0 9960 0 -1 -7769
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  sky130_fd_sc_hd__diode_2_2
timestamp 1715205430
transform 1 0 10144 0 -1 -7769
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  sky130_fd_sc_hd__diode_2_3
timestamp 1715205430
transform 1 0 10512 0 -1 -7769
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  sky130_fd_sc_hd__diode_2_4
timestamp 1715205430
transform 1 0 10696 0 -1 -7769
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1715205430
transform 1 0 9500 0 1 -8857
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1715205430
transform 1 0 9408 0 1 -8857
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1715205430
transform 1 0 10880 0 -1 -7769
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_2
timestamp 1715205430
transform 1 0 10880 0 1 -8857
box -38 -48 130 592
use sbvfcm  x1
timestamp 1719454670
transform 1 0 10300 0 1 -5200
box 5700 -4700 11200 5000
use output_amp  x2
timestamp 1719454661
transform 1 0 10400 0 -1 -14608
box 5100 -2900 11140 4900
use trim_res  x3
timestamp 1717344711
transform 1 0 8600 0 1 -15600
box 700 -3900 5534 -100
use sky130_fd_pr__nfet_01v8_2333C8  XM1
timestamp 1713045697
transform 1 0 11296 0 1 -5340
box -2196 -460 2196 460
use sky130_fd_pr__nfet_01v8_Q33MQV  XM2
timestamp 1717361709
transform 0 -1 14410 1 0 -6704
box -1196 -410 1196 410
use sky130_fd_pr__pfet_01v8_6H4ZLK  XM3
timestamp 1716081177
transform 0 1 13119 -1 0 -7204
box -1196 -719 1196 719
use sky130_fd_pr__pfet_01v8_B3G3L7  XM9
timestamp 1713056482
transform 0 -1 11837 1 0 -2475
box -2225 -2837 2225 2837
use sky130_fd_pr__pfet_01v8_XPMKX6  XM20
timestamp 1713045697
transform 0 1 9806 -1 0 -7352
box -226 -1219 226 1219
<< labels >>
rlabel via1 14900 -8000 15100 -7800 1 vref
rlabel via1 15800 -4200 16000 -4000 1 pbias
flabel metal1 21710 -10300 21910 -10100 0 FreeSans 256 0 0 0 vbg
port 0 nsew
flabel metal1 21710 -10600 21910 -10400 0 FreeSans 256 0 0 0 vbgtg
port 7 nsew
flabel metal1 21710 -10900 21910 -10700 0 FreeSans 256 0 0 0 vbgsc
port 6 nsew
flabel metal1 21710 -10000 21910 -9800 0 FreeSans 256 0 0 0 vptat
port 13 nsew
rlabel metal2 9360 -9330 9420 -9270 1 trim3buf
rlabel metal1 9360 -9390 9420 -9330 1 trim2buf
rlabel metal2 9360 -9450 9420 -9390 1 trim1buf
rlabel metal1 9360 -9510 9420 -9450 1 trim0buf
flabel metal1 8590 -8905 8790 -8705 0 FreeSans 256 0 0 0 dvss
port 4 nsew
flabel metal1 8590 -8600 8790 -8400 0 FreeSans 320 0 0 0 dvdd
port 14 nsew
rlabel metal1 8850 -7478 10806 -7434 1 avdd_ena
flabel metal1 8591 -7278 8791 -7078 0 FreeSans 256 0 0 0 avdd18
port 2 nsew
flabel metal1 8589 -8321 8788 -8121 0 FreeSans 256 0 0 0 ena
port 5 nsew
flabel metal1 8588 -8036 8788 -7836 0 FreeSans 256 0 0 0 trim3
port 8 nsew
flabel metal1 8589 -6570 8788 -6370 0 FreeSans 256 0 0 0 trim0
port 11 nsew
flabel metal1 8589 -6849 8788 -6649 0 FreeSans 256 0 0 0 trim1
port 10 nsew
flabel metal1 8589 -7763 8789 -7563 0 FreeSans 256 0 0 0 trim2
port 9 nsew
flabel metal1 21710 -11200 21910 -11000 0 FreeSans 256 0 0 0 avss
port 1 nsew
<< end >>
