magic
tech sky130A
magscale 1 2
timestamp 1713140876
<< pwell >>
rect -1756 -2472 1756 2472
<< psubdiff >>
rect -1720 2402 -1624 2436
rect 1624 2402 1720 2436
rect -1720 2340 -1686 2402
rect 1686 2340 1720 2402
rect -1720 -2402 -1686 -2340
rect 1686 -2402 1720 -2340
rect -1720 -2436 -1624 -2402
rect 1624 -2436 1720 -2402
<< psubdiffcont >>
rect -1624 2402 1624 2436
rect -1720 -2340 -1686 2340
rect 1686 -2340 1720 2340
rect -1624 -2436 1624 -2402
<< xpolycontact >>
rect -1590 1874 -1452 2306
rect -1590 -2306 -1452 -1874
rect -1356 1874 -1218 2306
rect -1356 -2306 -1218 -1874
rect -1122 1874 -984 2306
rect -1122 -2306 -984 -1874
rect -888 1874 -750 2306
rect -888 -2306 -750 -1874
rect -654 1874 -516 2306
rect -654 -2306 -516 -1874
rect -420 1874 -282 2306
rect -420 -2306 -282 -1874
rect -186 1874 -48 2306
rect -186 -2306 -48 -1874
rect 48 1874 186 2306
rect 48 -2306 186 -1874
rect 282 1874 420 2306
rect 282 -2306 420 -1874
rect 516 1874 654 2306
rect 516 -2306 654 -1874
rect 750 1874 888 2306
rect 750 -2306 888 -1874
rect 984 1874 1122 2306
rect 984 -2306 1122 -1874
rect 1218 1874 1356 2306
rect 1218 -2306 1356 -1874
rect 1452 1874 1590 2306
rect 1452 -2306 1590 -1874
<< xpolyres >>
rect -1590 -1874 -1452 1874
rect -1356 -1874 -1218 1874
rect -1122 -1874 -984 1874
rect -888 -1874 -750 1874
rect -654 -1874 -516 1874
rect -420 -1874 -282 1874
rect -186 -1874 -48 1874
rect 48 -1874 186 1874
rect 282 -1874 420 1874
rect 516 -1874 654 1874
rect 750 -1874 888 1874
rect 984 -1874 1122 1874
rect 1218 -1874 1356 1874
rect 1452 -1874 1590 1874
<< locali >>
rect -1720 2402 -1624 2436
rect 1624 2402 1720 2436
rect -1720 2340 -1686 2402
rect 1686 2340 1720 2402
rect -1720 -2402 -1686 -2340
rect 1686 -2402 1720 -2340
rect -1720 -2436 -1624 -2402
rect 1624 -2436 1720 -2402
<< viali >>
rect -1574 1891 -1468 2288
rect -1340 1891 -1234 2288
rect -1106 1891 -1000 2288
rect -872 1891 -766 2288
rect -638 1891 -532 2288
rect -404 1891 -298 2288
rect -170 1891 -64 2288
rect 64 1891 170 2288
rect 298 1891 404 2288
rect 532 1891 638 2288
rect 766 1891 872 2288
rect 1000 1891 1106 2288
rect 1234 1891 1340 2288
rect 1468 1891 1574 2288
rect -1574 -2288 -1468 -1891
rect -1340 -2288 -1234 -1891
rect -1106 -2288 -1000 -1891
rect -872 -2288 -766 -1891
rect -638 -2288 -532 -1891
rect -404 -2288 -298 -1891
rect -170 -2288 -64 -1891
rect 64 -2288 170 -1891
rect 298 -2288 404 -1891
rect 532 -2288 638 -1891
rect 766 -2288 872 -1891
rect 1000 -2288 1106 -1891
rect 1234 -2288 1340 -1891
rect 1468 -2288 1574 -1891
<< metal1 >>
rect -1580 2288 -1462 2300
rect -1580 1891 -1574 2288
rect -1468 1891 -1462 2288
rect -1580 1879 -1462 1891
rect -1346 2288 -1228 2300
rect -1346 1891 -1340 2288
rect -1234 1891 -1228 2288
rect -1346 1879 -1228 1891
rect -1112 2288 -994 2300
rect -1112 1891 -1106 2288
rect -1000 1891 -994 2288
rect -1112 1879 -994 1891
rect -878 2288 -760 2300
rect -878 1891 -872 2288
rect -766 1891 -760 2288
rect -878 1879 -760 1891
rect -644 2288 -526 2300
rect -644 1891 -638 2288
rect -532 1891 -526 2288
rect -644 1879 -526 1891
rect -410 2288 -292 2300
rect -410 1891 -404 2288
rect -298 1891 -292 2288
rect -410 1879 -292 1891
rect -176 2288 -58 2300
rect -176 1891 -170 2288
rect -64 1891 -58 2288
rect -176 1879 -58 1891
rect 58 2288 176 2300
rect 58 1891 64 2288
rect 170 1891 176 2288
rect 58 1879 176 1891
rect 292 2288 410 2300
rect 292 1891 298 2288
rect 404 1891 410 2288
rect 292 1879 410 1891
rect 526 2288 644 2300
rect 526 1891 532 2288
rect 638 1891 644 2288
rect 526 1879 644 1891
rect 760 2288 878 2300
rect 760 1891 766 2288
rect 872 1891 878 2288
rect 760 1879 878 1891
rect 994 2288 1112 2300
rect 994 1891 1000 2288
rect 1106 1891 1112 2288
rect 994 1879 1112 1891
rect 1228 2288 1346 2300
rect 1228 1891 1234 2288
rect 1340 1891 1346 2288
rect 1228 1879 1346 1891
rect 1462 2288 1580 2300
rect 1462 1891 1468 2288
rect 1574 1891 1580 2288
rect 1462 1879 1580 1891
rect -1580 -1891 -1462 -1879
rect -1580 -2288 -1574 -1891
rect -1468 -2288 -1462 -1891
rect -1580 -2300 -1462 -2288
rect -1346 -1891 -1228 -1879
rect -1346 -2288 -1340 -1891
rect -1234 -2288 -1228 -1891
rect -1346 -2300 -1228 -2288
rect -1112 -1891 -994 -1879
rect -1112 -2288 -1106 -1891
rect -1000 -2288 -994 -1891
rect -1112 -2300 -994 -2288
rect -878 -1891 -760 -1879
rect -878 -2288 -872 -1891
rect -766 -2288 -760 -1891
rect -878 -2300 -760 -2288
rect -644 -1891 -526 -1879
rect -644 -2288 -638 -1891
rect -532 -2288 -526 -1891
rect -644 -2300 -526 -2288
rect -410 -1891 -292 -1879
rect -410 -2288 -404 -1891
rect -298 -2288 -292 -1891
rect -410 -2300 -292 -2288
rect -176 -1891 -58 -1879
rect -176 -2288 -170 -1891
rect -64 -2288 -58 -1891
rect -176 -2300 -58 -2288
rect 58 -1891 176 -1879
rect 58 -2288 64 -1891
rect 170 -2288 176 -1891
rect 58 -2300 176 -2288
rect 292 -1891 410 -1879
rect 292 -2288 298 -1891
rect 404 -2288 410 -1891
rect 292 -2300 410 -2288
rect 526 -1891 644 -1879
rect 526 -2288 532 -1891
rect 638 -2288 644 -1891
rect 526 -2300 644 -2288
rect 760 -1891 878 -1879
rect 760 -2288 766 -1891
rect 872 -2288 878 -1891
rect 760 -2300 878 -2288
rect 994 -1891 1112 -1879
rect 994 -2288 1000 -1891
rect 1106 -2288 1112 -1891
rect 994 -2300 1112 -2288
rect 1228 -1891 1346 -1879
rect 1228 -2288 1234 -1891
rect 1340 -2288 1346 -1891
rect 1228 -2300 1346 -2288
rect 1462 -1891 1580 -1879
rect 1462 -2288 1468 -1891
rect 1574 -2288 1580 -1891
rect 1462 -2300 1580 -2288
<< properties >>
string FIXED_BBOX -1703 -2419 1703 2419
string gencell sky130_fd_pr__res_xhigh_po_0p69
string library sky130
string parameters w 0.690 l 18.9 m 1 nx 14 wmin 0.690 lmin 0.50 rho 2000 val 55.328k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.690 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
