magic
tech sky130A
magscale 1 2
timestamp 1713049709
<< nwell >>
rect -1225 -4219 1225 4219
<< pmos >>
rect -1029 -4000 -29 4000
rect 29 -4000 1029 4000
<< pdiff >>
rect -1087 3988 -1029 4000
rect -1087 -3988 -1075 3988
rect -1041 -3988 -1029 3988
rect -1087 -4000 -1029 -3988
rect -29 3988 29 4000
rect -29 -3988 -17 3988
rect 17 -3988 29 3988
rect -29 -4000 29 -3988
rect 1029 3988 1087 4000
rect 1029 -3988 1041 3988
rect 1075 -3988 1087 3988
rect 1029 -4000 1087 -3988
<< pdiffc >>
rect -1075 -3988 -1041 3988
rect -17 -3988 17 3988
rect 1041 -3988 1075 3988
<< nsubdiff >>
rect -1189 4149 -1093 4183
rect 1093 4149 1189 4183
rect -1189 4087 -1155 4149
rect 1155 4087 1189 4149
rect -1189 -4149 -1155 -4087
rect 1155 -4149 1189 -4087
rect -1189 -4183 -1093 -4149
rect 1093 -4183 1189 -4149
<< nsubdiffcont >>
rect -1093 4149 1093 4183
rect -1189 -4087 -1155 4087
rect 1155 -4087 1189 4087
rect -1093 -4183 1093 -4149
<< poly >>
rect -1029 4081 -29 4097
rect -1029 4047 -1013 4081
rect -45 4047 -29 4081
rect -1029 4000 -29 4047
rect 29 4081 1029 4097
rect 29 4047 45 4081
rect 1013 4047 1029 4081
rect 29 4000 1029 4047
rect -1029 -4047 -29 -4000
rect -1029 -4081 -1013 -4047
rect -45 -4081 -29 -4047
rect -1029 -4097 -29 -4081
rect 29 -4047 1029 -4000
rect 29 -4081 45 -4047
rect 1013 -4081 1029 -4047
rect 29 -4097 1029 -4081
<< polycont >>
rect -1013 4047 -45 4081
rect 45 4047 1013 4081
rect -1013 -4081 -45 -4047
rect 45 -4081 1013 -4047
<< locali >>
rect -1189 4149 -1093 4183
rect 1093 4149 1189 4183
rect -1189 4087 -1155 4149
rect 1155 4087 1189 4149
rect -1029 4047 -1013 4081
rect -45 4047 -29 4081
rect 29 4047 45 4081
rect 1013 4047 1029 4081
rect -1075 3988 -1041 4004
rect -1075 -4004 -1041 -3988
rect -17 3988 17 4004
rect -17 -4004 17 -3988
rect 1041 3988 1075 4004
rect 1041 -4004 1075 -3988
rect -1029 -4081 -1013 -4047
rect -45 -4081 -29 -4047
rect 29 -4081 45 -4047
rect 1013 -4081 1029 -4047
rect -1189 -4149 -1155 -4087
rect 1155 -4149 1189 -4087
rect -1189 -4183 -1093 -4149
rect 1093 -4183 1189 -4149
<< viali >>
rect -1013 4047 -45 4081
rect 45 4047 1013 4081
rect -1075 -3988 -1041 3988
rect -17 -3988 17 3988
rect 1041 -3988 1075 3988
rect -1013 -4081 -45 -4047
rect 45 -4081 1013 -4047
<< metal1 >>
rect -1025 4081 -33 4087
rect -1025 4047 -1013 4081
rect -45 4047 -33 4081
rect -1025 4041 -33 4047
rect 33 4081 1025 4087
rect 33 4047 45 4081
rect 1013 4047 1025 4081
rect 33 4041 1025 4047
rect -1081 3988 -1035 4000
rect -1081 -3988 -1075 3988
rect -1041 -3988 -1035 3988
rect -1081 -4000 -1035 -3988
rect -23 3988 23 4000
rect -23 -3988 -17 3988
rect 17 -3988 23 3988
rect -23 -4000 23 -3988
rect 1035 3988 1081 4000
rect 1035 -3988 1041 3988
rect 1075 -3988 1081 3988
rect 1035 -4000 1081 -3988
rect -1025 -4047 -33 -4041
rect -1025 -4081 -1013 -4047
rect -45 -4081 -33 -4047
rect -1025 -4087 -33 -4081
rect 33 -4047 1025 -4041
rect 33 -4081 45 -4047
rect 1013 -4081 1025 -4047
rect 33 -4087 1025 -4081
<< properties >>
string FIXED_BBOX -1172 -4166 1172 4166
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 40.0 l 5.0 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
