magic
tech sky130A
magscale 1 2
timestamp 1713051387
<< pwell >>
rect -235 -1272 235 1272
<< psubdiff >>
rect -199 1202 -103 1236
rect 103 1202 199 1236
rect -199 1140 -165 1202
rect 165 1140 199 1202
rect -199 -1202 -165 -1140
rect 165 -1202 199 -1140
rect -199 -1236 -103 -1202
rect 103 -1236 199 -1202
<< psubdiffcont >>
rect -103 1202 103 1236
rect -199 -1140 -165 1140
rect 165 -1140 199 1140
rect -103 -1236 103 -1202
<< xpolycontact >>
rect -69 674 69 1106
rect -69 -1106 69 -674
<< xpolyres >>
rect -69 -674 69 674
<< locali >>
rect -199 1202 -103 1236
rect 103 1202 199 1236
rect -199 1140 -165 1202
rect 165 1140 199 1202
rect -199 -1202 -165 -1140
rect 165 -1202 199 -1140
rect -199 -1236 -103 -1202
rect 103 -1236 199 -1202
<< viali >>
rect -53 691 53 1088
rect -53 -1088 53 -691
<< metal1 >>
rect -59 1088 59 1100
rect -59 691 -53 1088
rect 53 691 59 1088
rect -59 679 59 691
rect -59 -691 59 -679
rect -59 -1088 -53 -691
rect 53 -1088 59 -691
rect -59 -1100 59 -1088
<< properties >>
string FIXED_BBOX -182 -1219 182 1219
string gencell sky130_fd_pr__res_xhigh_po_0p69
string library sky130
string parameters w 0.690 l 6.9 m 1 nx 1 wmin 0.690 lmin 0.50 rho 2000 val 20.545k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.690 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
