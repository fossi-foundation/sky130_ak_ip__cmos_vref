magic
tech sky130A
magscale 1 2
timestamp 1713146894
<< error_p >>
rect 20500 -14708 20506 -14702
rect 20694 -14708 20700 -14702
rect 20494 -14714 20500 -14708
rect 20700 -14714 20706 -14708
rect 20494 -14908 20500 -14902
rect 20500 -14914 20506 -14908
<< error_s >>
rect 15597 -1200 15655 -1194
rect 15597 -1234 15609 -1200
rect 15597 -1240 15655 -1234
rect 16100 -1564 16106 -808
rect 15597 -3328 15655 -3322
rect 15597 -3362 15609 -3328
rect 15597 -3368 15655 -3362
rect 14600 -8600 14606 -8594
rect 14594 -8606 14600 -8600
rect 14594 -8800 14600 -8794
rect 14600 -8806 14606 -8800
rect 19600 -9500 19606 -9494
rect 19794 -9500 19800 -9494
rect 19594 -9506 19600 -9500
rect 19800 -9506 19806 -9500
rect 19800 -9700 19806 -9694
rect 19794 -9706 19800 -9700
rect 17900 -10400 17906 -10394
rect 18094 -10400 18100 -10394
rect 17894 -10406 17900 -10400
rect 18100 -10406 18106 -10400
rect 14900 -11700 14906 -11694
rect 15094 -11700 15100 -11694
rect 14894 -11706 14900 -11700
rect 15100 -11706 15106 -11700
rect 19600 -11708 19606 -11702
rect 19794 -11708 19800 -11702
rect 19594 -11714 19600 -11708
rect 19800 -11714 19806 -11708
rect 14894 -11900 14900 -11894
rect 15100 -11900 15106 -11894
rect 14900 -11906 14906 -11900
rect 15094 -11906 15100 -11900
rect 19594 -11908 19600 -11902
rect 19800 -11908 19806 -11902
rect 19600 -11914 19606 -11908
rect 19794 -11914 19800 -11908
rect 17500 -12008 17506 -12002
rect 17694 -12008 17700 -12002
rect 17494 -12014 17500 -12008
rect 17700 -12014 17706 -12008
rect 17494 -12208 17500 -12202
rect 17700 -12208 17706 -12202
rect 17500 -12214 17506 -12208
rect 17694 -12214 17700 -12208
rect 19000 -13408 19006 -13402
rect 19194 -13408 19200 -13402
rect 18994 -13414 19000 -13408
rect 19200 -13414 19206 -13408
rect 18994 -13608 19000 -13602
rect 19200 -13608 19206 -13602
rect 19000 -13614 19006 -13608
rect 19194 -13614 19200 -13608
rect 10980 -16246 10986 -16240
rect 11174 -16246 11180 -16240
rect 10974 -16252 10980 -16246
rect 11180 -16252 11186 -16246
rect 10974 -16446 10980 -16440
rect 11180 -16446 11186 -16440
rect 10980 -16452 10986 -16446
rect 11174 -16452 11180 -16446
rect 14140 -16560 14146 -16554
rect 14334 -16560 14340 -16554
rect 14134 -16566 14140 -16560
rect 14340 -16566 14346 -16560
rect 13140 -16592 13146 -16586
rect 13146 -16598 13152 -16592
rect 14134 -16760 14140 -16755
rect 14340 -16760 14346 -16755
rect 14140 -16766 14146 -16760
rect 14334 -16766 14340 -16760
<< metal1 >>
rect 15500 -900 15700 -700
rect 15800 -900 16000 -700
rect 9000 -8500 9200 -8300
rect 15800 -8600 16000 -6900
rect 9000 -8800 9200 -8600
rect 14800 -8800 16000 -8600
rect 9000 -9100 14300 -8900
rect 14500 -9100 16000 -8900
rect 13500 -9500 14800 -9300
rect 13500 -10000 14500 -9800
rect 13600 -10500 14200 -10300
rect 14000 -10700 14200 -10500
rect 14300 -10400 14500 -10000
rect 14600 -10100 14800 -9500
rect 15800 -9500 16000 -9100
rect 19194 -9200 19200 -9000
rect 19400 -9200 19406 -9000
rect 19520 -9500 19720 -9054
rect 15800 -9700 19600 -9500
rect 17100 -10000 18700 -9800
rect 18900 -10000 18906 -9800
rect 14600 -10300 21500 -10100
rect 14300 -10600 17900 -10400
rect 18100 -10600 21500 -10400
rect 14000 -10900 21500 -10700
rect 15800 -11400 16000 -10900
rect 19200 -11000 19400 -10994
rect 19400 -11200 21500 -11000
rect 19200 -11206 19400 -11200
rect 13600 -11600 15400 -11400
rect 17894 -11500 17900 -11300
rect 18100 -11500 18106 -11300
rect 14300 -11700 14500 -11694
rect 11640 -14700 13400 -14500
rect 11640 -15060 11840 -14700
rect 14300 -14860 14500 -11900
rect 11900 -15060 14500 -14860
rect 14600 -11700 14800 -11694
rect 9000 -15300 9200 -15100
rect 9000 -15600 9200 -15400
rect 14600 -16608 14800 -11900
rect 14900 -16308 15100 -11900
rect 15200 -16008 15400 -11600
rect 18700 -11708 18900 -11702
rect 18700 -11914 18900 -11908
rect 15200 -16208 15700 -16008
rect 14900 -16508 15700 -16308
rect 14600 -16808 15700 -16608
rect 9000 -19200 9200 -19000
rect 9000 -19500 9200 -19300
<< via1 >>
rect 14600 -8800 14800 -8600
rect 14300 -9100 14500 -8900
rect 19200 -9200 19400 -9000
rect 19600 -9700 19800 -9500
rect 18700 -10000 18900 -9800
rect 17900 -10600 18100 -10400
rect 19200 -11200 19400 -11000
rect 17900 -11500 18100 -11300
rect 14300 -11900 14500 -11700
rect 14600 -11900 14800 -11700
rect 14900 -11900 15100 -11700
rect 18700 -11908 18900 -11708
rect 19600 -11908 19800 -11708
<< metal2 >>
rect 14600 -8600 14800 -8500
rect 14300 -8900 14500 -8893
rect 14300 -11700 14500 -9100
rect 14600 -11700 14800 -8800
rect 14900 -11700 15100 -8500
rect 19200 -9000 19400 -8994
rect 18700 -9800 18900 -9794
rect 17900 -11300 18100 -10600
rect 17900 -11506 18100 -11500
rect 14294 -11900 14300 -11700
rect 14500 -11900 14506 -11700
rect 14594 -11900 14600 -11700
rect 14800 -11900 14806 -11700
rect 18700 -11708 18900 -10000
rect 19200 -11000 19400 -9200
rect 19194 -11200 19200 -11000
rect 19400 -11200 19406 -11000
rect 19600 -11708 19800 -9700
rect 18694 -11908 18700 -11708
rect 18900 -11908 18906 -11708
use sky130_fd_pr__res_xhigh_po_0p69_E9MCU4  R1
timestamp 1713140876
transform 0 1 11399 -1 0 -9631
box -469 -2399 469 2399
use sky130_fd_pr__res_xhigh_po_0p69_39QBTQ  R2
timestamp 1713056482
transform 0 1 16942 -1 0 -11365
box -235 -1442 235 1442
use sky130_fd_pr__res_xhigh_po_0p69_NB3ZKH  R3
timestamp 1713140876
transform 0 1 11445 -1 0 -10714
box -586 -2445 586 2445
use sky130_fd_pr__res_xhigh_po_0p69_GAZAU4  R4
timestamp 1713140876
transform 0 -1 11472 1 0 -13044
box -1756 -2472 1756 2472
use sbvfcm  x1
timestamp 1713048788
transform 1 0 10398 0 1 -5204
box 5702 -4196 11000 5078
use output_amp  x2
timestamp 1713128983
transform 1 0 10400 0 -1 -14608
box 5100 -2903 11100 4892
use trim_res  x3
timestamp 1713116496
transform 1 0 8480 0 1 -15320
box 720 -4180 5972 460
use sky130_fd_pr__nfet_01v8_2333C8  XM1
timestamp 1713045697
transform 1 0 11196 0 1 -7540
box -2196 -460 2196 460
use sky130_fd_pr__nfet_01v8_QXBCRM  XM2
timestamp 1713051622
transform 1 0 10196 0 1 -6690
box -1196 -310 1196 310
use sky130_fd_pr__pfet_01v8_6H4ZLK  XM3
timestamp 1713045697
transform 0 1 14219 -1 0 -6804
box -1196 -719 1196 719
use sky130_fd_pr__pfet_01v8_B3G3L7  XM9
timestamp 1713056482
transform 0 -1 11937 1 0 -3075
box -2225 -2837 2225 2837
use sky130_fd_pr__pfet_01v8_XPMKX6  XM20
timestamp 1713045697
transform 1 0 15626 0 1 -2281
box -226 -1219 226 1219
<< labels >>
flabel metal1 21300 -10300 21500 -10100 0 FreeSans 256 0 0 0 vbg
port 0 nsew
flabel metal1 21300 -10600 21500 -10400 0 FreeSans 256 0 0 0 vbgtg
port 7 nsew
flabel metal1 21300 -10900 21500 -10700 0 FreeSans 256 0 0 0 vbgsc
port 6 nsew
flabel metal1 15800 -900 16000 -700 0 FreeSans 256 0 0 0 avdd18
port 2 nsew
flabel metal1 15500 -900 15700 -700 0 FreeSans 256 0 0 0 ena
port 5 nsew
flabel metal1 21300 -11200 21500 -11000 0 FreeSans 256 0 0 0 vptat
port 13 nsew
flabel metal1 9000 -19500 9200 -19300 0 FreeSans 256 0 0 0 trim3
port 8 nsew
flabel metal1 9000 -19200 9200 -19000 0 FreeSans 256 0 0 0 trim2
port 9 nsew
flabel metal1 9000 -15600 9200 -15400 0 FreeSans 256 0 0 0 trim0
port 11 nsew
flabel metal1 9000 -15300 9200 -15100 0 FreeSans 256 0 0 0 trim1
port 10 nsew
flabel metal1 9000 -9100 9200 -8900 0 FreeSans 256 0 0 0 avss
port 1 nsew
flabel metal1 9000 -8800 9200 -8600 0 FreeSans 256 0 0 0 dvss
port 4 nsew
flabel metal1 9000 -8500 9200 -8300 0 FreeSans 256 0 0 0 dvdd
port 3 nsew
<< end >>
