magic
tech sky130A
magscale 1 2
timestamp 1713214705
<< error_s >>
rect 5972 4100 6000 4106
rect 10900 4100 10920 4106
rect 6000 4072 6028 4078
rect 10872 4072 10892 4078
rect 6900 3500 6906 3506
rect 6894 3494 6900 3500
rect 6894 3300 6900 3306
rect 7100 3300 7106 3306
rect 6900 3294 6906 3300
rect 7094 3294 7100 3300
rect 6900 2200 6906 2206
rect 6894 2194 6900 2200
rect 6894 2000 6900 2006
rect 6900 1994 6906 2000
rect 10874 1194 10900 1406
rect 10902 1166 10928 1434
rect 8000 1000 8020 1006
rect 8872 1000 8900 1006
rect 7972 972 7992 978
rect 8900 972 8928 978
rect 8800 600 8806 606
rect 8994 600 9000 606
rect 8794 594 8800 600
rect 9000 594 9006 600
rect 8794 400 8800 406
rect 9000 400 9006 406
rect 8800 394 8806 400
rect 8994 394 9000 400
rect 8700 100 8706 106
rect 8894 100 8900 106
rect 8694 94 8700 100
rect 8900 94 8906 100
rect 8694 -100 8700 -94
rect 8700 -106 8706 -100
rect 9072 -500 9100 -494
rect 9100 -528 9128 -522
rect 7700 -1000 7706 -994
rect 7894 -1000 7900 -994
rect 7694 -1006 7700 -1000
rect 7900 -1006 7906 -1000
rect 7694 -1200 7700 -1194
rect 7900 -1200 7906 -1194
rect 7700 -1206 7706 -1200
rect 7894 -1206 7900 -1200
rect 7700 -2000 7706 -1994
rect 7894 -2000 7900 -1994
rect 7694 -2006 7700 -2000
rect 7900 -2006 7906 -2000
rect 7694 -2200 7700 -2194
rect 7900 -2200 7906 -2194
rect 7700 -2206 7706 -2200
rect 7894 -2206 7900 -2200
<< metal1 >>
rect 5700 5300 11200 5500
rect 5700 5100 5900 5300
rect 5700 4100 6000 5100
rect 6900 4700 7100 5200
rect 6900 4500 8400 4700
rect 5700 3600 5900 4100
rect 6900 3500 7100 4500
rect 5700 3300 6900 3500
rect 6900 2200 7100 3100
rect 8200 3000 8400 4500
rect 5900 1200 6000 1400
rect 6200 1200 6206 1400
rect 6900 700 7100 2000
rect 8000 1000 8400 3000
rect 8500 4500 8900 4700
rect 8500 3000 8700 4500
rect 9800 3500 10000 5200
rect 11000 5100 11200 5300
rect 10900 4100 11200 5100
rect 9800 3294 10000 3300
rect 8500 1000 8900 3000
rect 9800 2200 10000 3100
rect 9800 900 10000 2000
rect 10700 1400 10900 1406
rect 10700 1194 10900 1200
rect 5700 500 7100 700
rect 6094 200 6100 400
rect 6300 200 6306 400
rect 5700 -100 8700 100
rect 5700 -3400 5900 -100
rect 7694 -400 7700 -200
rect 7900 -400 7906 -200
rect 6100 -600 6300 -594
rect 6100 -806 6300 -800
rect 6094 -1700 6100 -1500
rect 6300 -1700 6306 -1500
rect 6094 -2600 6100 -2400
rect 6300 -2600 6306 -2400
rect 7694 -3100 7700 -2900
rect 7900 -3100 7906 -2900
rect 8700 -3300 8900 -100
rect 9000 -500 9100 500
rect 9200 100 9400 600
rect 9600 400 9700 500
rect 9200 -600 9400 -100
rect 9500 -400 9700 400
rect 9600 -800 9700 -400
rect 9300 -1000 9700 -800
rect 6100 -3500 6300 -3300
rect 6094 -3700 6100 -3500
rect 6300 -3700 9200 -3500
rect 9300 -3700 9500 -1000
rect 11000 -2900 11200 4100
<< via1 >>
rect 6900 3300 7100 3500
rect 6900 2000 7100 2200
rect 6000 1200 6200 1400
rect 9800 3300 10000 3500
rect 9800 2000 10000 2200
rect 10700 1200 10900 1400
rect 8800 400 9000 600
rect 6100 200 6300 400
rect 8700 -100 8900 100
rect 7700 -400 7900 -200
rect 6100 -800 6300 -600
rect 7700 -1200 7900 -1000
rect 6100 -1700 6300 -1500
rect 7700 -2200 7900 -2000
rect 6100 -2600 6300 -2400
rect 7700 -3100 7900 -2900
rect 9200 -100 9400 100
rect 6100 -3700 6300 -3500
<< metal2 >>
rect 7100 3300 9800 3500
rect 10000 3300 10006 3500
rect 7100 2000 9800 2200
rect 10000 2000 10006 2200
rect 6000 1400 6200 1406
rect 6200 1200 7900 1400
rect 6000 1194 6200 1200
rect 6100 400 6300 406
rect 6100 -600 6300 200
rect 7700 -200 7900 1200
rect 8800 1200 10700 1400
rect 10900 1200 10906 1400
rect 8800 600 9000 1200
rect 8900 -100 9200 100
rect 9400 -100 9406 100
rect 6094 -800 6100 -600
rect 6300 -800 6306 -600
rect 6100 -1500 6300 -800
rect 6100 -2400 6300 -1700
rect 6100 -3500 6300 -2600
rect 7700 -1000 7900 -400
rect 7700 -2000 7900 -1200
rect 7700 -2900 7900 -2200
rect 7700 -3106 7900 -3100
rect 6100 -3706 6300 -3700
use sky130_fd_pr__nfet_01v8_QTPFY2  sky130_fd_pr__nfet_01v8_QTPFY2_0
timestamp 1713212409
transform 0 1 7260 -1 0 -1601
box -1999 -1460 1999 1460
use sky130_fd_pr__cap_mim_m3_1_VCAG9S  XC1
timestamp 1713045697
transform -1 0 10386 0 -1 -2760
box -686 -540 686 540
use sky130_fd_pr__nfet_01v8_QGRVRG  XM4
timestamp 1713045697
transform 1 0 9296 0 1 10
box -396 -710 396 710
use sky130_fd_pr__nfet_01v8_ME6MQD  XM5
timestamp 1713045697
transform 1 0 6996 0 1 2010
box -1196 -1210 1196 1210
use sky130_fd_pr__nfet_01v8_ME6MQD  XM6
timestamp 1713045697
transform 1 0 9896 0 1 2010
box -1196 -1210 1196 1210
use sky130_fd_pr__pfet_01v8_6H4ZLK  XM7
timestamp 1713045697
transform 1 0 6996 0 1 4619
box -1196 -719 1196 719
use sky130_fd_pr__pfet_01v8_6H4ZLK  XM8
timestamp 1713045697
transform 1 0 9896 0 1 4619
box -1196 -719 1196 719
use sky130_fd_pr__nfet_01v8_TTEWAE  XM10
timestamp 1713212409
transform 1 0 10396 0 1 10
box -696 -710 696 710
use sky130_fd_pr__nfet_01v8_BSH2JQ  XM11
timestamp 1713212409
transform -1 0 10396 0 -1 -1490
box -696 -710 696 710
<< labels >>
flabel metal1 5700 3300 5900 3500 0 FreeSans 256 0 0 0 pbias
port 1 nsew
flabel metal1 5700 3600 5900 3800 0 FreeSans 256 0 0 0 vdd
port 0 nsew
flabel metal1 5700 500 5900 700 0 FreeSans 256 0 0 0 nbias
port 2 nsew
flabel metal1 9000 -3700 9200 -3500 0 FreeSans 256 0 0 0 vx
port 3 nsew
flabel metal1 9300 -3700 9500 -3500 0 FreeSans 256 0 0 0 vss
port 4 nsew
<< end >>
