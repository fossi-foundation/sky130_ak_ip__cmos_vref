magic
tech sky130A
magscale 1 2
timestamp 1713049709
<< nwell >>
rect -696 -8337 696 8337
<< pmos >>
rect -500 118 500 8118
rect -500 -8118 500 -118
<< pdiff >>
rect -558 8106 -500 8118
rect -558 130 -546 8106
rect -512 130 -500 8106
rect -558 118 -500 130
rect 500 8106 558 8118
rect 500 130 512 8106
rect 546 130 558 8106
rect 500 118 558 130
rect -558 -130 -500 -118
rect -558 -8106 -546 -130
rect -512 -8106 -500 -130
rect -558 -8118 -500 -8106
rect 500 -130 558 -118
rect 500 -8106 512 -130
rect 546 -8106 558 -130
rect 500 -8118 558 -8106
<< pdiffc >>
rect -546 130 -512 8106
rect 512 130 546 8106
rect -546 -8106 -512 -130
rect 512 -8106 546 -130
<< nsubdiff >>
rect -660 8267 -564 8301
rect 564 8267 660 8301
rect -660 8205 -626 8267
rect 626 8205 660 8267
rect -660 -8267 -626 -8205
rect 626 -8267 660 -8205
rect -660 -8301 -564 -8267
rect 564 -8301 660 -8267
<< nsubdiffcont >>
rect -564 8267 564 8301
rect -660 -8205 -626 8205
rect 626 -8205 660 8205
rect -564 -8301 564 -8267
<< poly >>
rect -500 8199 500 8215
rect -500 8165 -484 8199
rect 484 8165 500 8199
rect -500 8118 500 8165
rect -500 71 500 118
rect -500 37 -484 71
rect 484 37 500 71
rect -500 21 500 37
rect -500 -37 500 -21
rect -500 -71 -484 -37
rect 484 -71 500 -37
rect -500 -118 500 -71
rect -500 -8165 500 -8118
rect -500 -8199 -484 -8165
rect 484 -8199 500 -8165
rect -500 -8215 500 -8199
<< polycont >>
rect -484 8165 484 8199
rect -484 37 484 71
rect -484 -71 484 -37
rect -484 -8199 484 -8165
<< locali >>
rect -660 8267 -564 8301
rect 564 8267 660 8301
rect -660 8205 -626 8267
rect 626 8205 660 8267
rect -500 8165 -484 8199
rect 484 8165 500 8199
rect -546 8106 -512 8122
rect -546 114 -512 130
rect 512 8106 546 8122
rect 512 114 546 130
rect -500 37 -484 71
rect 484 37 500 71
rect -500 -71 -484 -37
rect 484 -71 500 -37
rect -546 -130 -512 -114
rect -546 -8122 -512 -8106
rect 512 -130 546 -114
rect 512 -8122 546 -8106
rect -500 -8199 -484 -8165
rect 484 -8199 500 -8165
rect -660 -8267 -626 -8205
rect 626 -8267 660 -8205
rect -660 -8301 -564 -8267
rect 564 -8301 660 -8267
<< viali >>
rect -484 8165 484 8199
rect -546 130 -512 8106
rect 512 130 546 8106
rect -484 37 484 71
rect -484 -71 484 -37
rect -546 -8106 -512 -130
rect 512 -8106 546 -130
rect -484 -8199 484 -8165
<< metal1 >>
rect -496 8199 496 8205
rect -496 8165 -484 8199
rect 484 8165 496 8199
rect -496 8159 496 8165
rect -552 8106 -506 8118
rect -552 130 -546 8106
rect -512 130 -506 8106
rect -552 118 -506 130
rect 506 8106 552 8118
rect 506 130 512 8106
rect 546 130 552 8106
rect 506 118 552 130
rect -496 71 496 77
rect -496 37 -484 71
rect 484 37 496 71
rect -496 31 496 37
rect -496 -37 496 -31
rect -496 -71 -484 -37
rect 484 -71 496 -37
rect -496 -77 496 -71
rect -552 -130 -506 -118
rect -552 -8106 -546 -130
rect -512 -8106 -506 -130
rect -552 -8118 -506 -8106
rect 506 -130 552 -118
rect 506 -8106 512 -130
rect 546 -8106 552 -130
rect 506 -8118 552 -8106
rect -496 -8165 496 -8159
rect -496 -8199 -484 -8165
rect 484 -8199 496 -8165
rect -496 -8205 496 -8199
<< properties >>
string FIXED_BBOX -643 -8284 643 8284
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 40.0 l 5.0 m 2 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
