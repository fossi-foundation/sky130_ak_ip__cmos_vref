magic
tech sky130A
magscale 1 2
timestamp 1713052702
<< nwell >>
rect -2225 -2337 2225 2337
<< pmos >>
rect -2029 118 -29 2118
rect 29 118 2029 2118
rect -2029 -2118 -29 -118
rect 29 -2118 2029 -118
<< pdiff >>
rect -2087 2106 -2029 2118
rect -2087 130 -2075 2106
rect -2041 130 -2029 2106
rect -2087 118 -2029 130
rect -29 2106 29 2118
rect -29 130 -17 2106
rect 17 130 29 2106
rect -29 118 29 130
rect 2029 2106 2087 2118
rect 2029 130 2041 2106
rect 2075 130 2087 2106
rect 2029 118 2087 130
rect -2087 -130 -2029 -118
rect -2087 -2106 -2075 -130
rect -2041 -2106 -2029 -130
rect -2087 -2118 -2029 -2106
rect -29 -130 29 -118
rect -29 -2106 -17 -130
rect 17 -2106 29 -130
rect -29 -2118 29 -2106
rect 2029 -130 2087 -118
rect 2029 -2106 2041 -130
rect 2075 -2106 2087 -130
rect 2029 -2118 2087 -2106
<< pdiffc >>
rect -2075 130 -2041 2106
rect -17 130 17 2106
rect 2041 130 2075 2106
rect -2075 -2106 -2041 -130
rect -17 -2106 17 -130
rect 2041 -2106 2075 -130
<< nsubdiff >>
rect -2189 2267 -2093 2301
rect 2093 2267 2189 2301
rect -2189 2205 -2155 2267
rect 2155 2205 2189 2267
rect -2189 -2267 -2155 -2205
rect 2155 -2267 2189 -2205
rect -2189 -2301 -2093 -2267
rect 2093 -2301 2189 -2267
<< nsubdiffcont >>
rect -2093 2267 2093 2301
rect -2189 -2205 -2155 2205
rect 2155 -2205 2189 2205
rect -2093 -2301 2093 -2267
<< poly >>
rect -2029 2199 -29 2215
rect -2029 2165 -2013 2199
rect -45 2165 -29 2199
rect -2029 2118 -29 2165
rect 29 2199 2029 2215
rect 29 2165 45 2199
rect 2013 2165 2029 2199
rect 29 2118 2029 2165
rect -2029 71 -29 118
rect -2029 37 -2013 71
rect -45 37 -29 71
rect -2029 21 -29 37
rect 29 71 2029 118
rect 29 37 45 71
rect 2013 37 2029 71
rect 29 21 2029 37
rect -2029 -37 -29 -21
rect -2029 -71 -2013 -37
rect -45 -71 -29 -37
rect -2029 -118 -29 -71
rect 29 -37 2029 -21
rect 29 -71 45 -37
rect 2013 -71 2029 -37
rect 29 -118 2029 -71
rect -2029 -2165 -29 -2118
rect -2029 -2199 -2013 -2165
rect -45 -2199 -29 -2165
rect -2029 -2215 -29 -2199
rect 29 -2165 2029 -2118
rect 29 -2199 45 -2165
rect 2013 -2199 2029 -2165
rect 29 -2215 2029 -2199
<< polycont >>
rect -2013 2165 -45 2199
rect 45 2165 2013 2199
rect -2013 37 -45 71
rect 45 37 2013 71
rect -2013 -71 -45 -37
rect 45 -71 2013 -37
rect -2013 -2199 -45 -2165
rect 45 -2199 2013 -2165
<< locali >>
rect -2189 2267 -2093 2301
rect 2093 2267 2189 2301
rect -2189 2205 -2155 2267
rect 2155 2205 2189 2267
rect -2029 2165 -2013 2199
rect -45 2165 -29 2199
rect 29 2165 45 2199
rect 2013 2165 2029 2199
rect -2075 2106 -2041 2122
rect -2075 114 -2041 130
rect -17 2106 17 2122
rect -17 114 17 130
rect 2041 2106 2075 2122
rect 2041 114 2075 130
rect -2029 37 -2013 71
rect -45 37 -29 71
rect 29 37 45 71
rect 2013 37 2029 71
rect -2029 -71 -2013 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 2013 -71 2029 -37
rect -2075 -130 -2041 -114
rect -2075 -2122 -2041 -2106
rect -17 -130 17 -114
rect -17 -2122 17 -2106
rect 2041 -130 2075 -114
rect 2041 -2122 2075 -2106
rect -2029 -2199 -2013 -2165
rect -45 -2199 -29 -2165
rect 29 -2199 45 -2165
rect 2013 -2199 2029 -2165
rect -2189 -2267 -2155 -2205
rect 2155 -2267 2189 -2205
rect -2189 -2301 -2093 -2267
rect 2093 -2301 2189 -2267
<< viali >>
rect -2013 2165 -45 2199
rect 45 2165 2013 2199
rect -2075 130 -2041 2106
rect -17 130 17 2106
rect 2041 130 2075 2106
rect -2013 37 -45 71
rect 45 37 2013 71
rect -2013 -71 -45 -37
rect 45 -71 2013 -37
rect -2075 -2106 -2041 -130
rect -17 -2106 17 -130
rect 2041 -2106 2075 -130
rect -2013 -2199 -45 -2165
rect 45 -2199 2013 -2165
<< metal1 >>
rect -2025 2199 -33 2205
rect -2025 2165 -2013 2199
rect -45 2165 -33 2199
rect -2025 2159 -33 2165
rect 33 2199 2025 2205
rect 33 2165 45 2199
rect 2013 2165 2025 2199
rect 33 2159 2025 2165
rect -2081 2106 -2035 2118
rect -2081 130 -2075 2106
rect -2041 130 -2035 2106
rect -2081 118 -2035 130
rect -23 2106 23 2118
rect -23 130 -17 2106
rect 17 130 23 2106
rect -23 118 23 130
rect 2035 2106 2081 2118
rect 2035 130 2041 2106
rect 2075 130 2081 2106
rect 2035 118 2081 130
rect -2025 71 -33 77
rect -2025 37 -2013 71
rect -45 37 -33 71
rect -2025 31 -33 37
rect 33 71 2025 77
rect 33 37 45 71
rect 2013 37 2025 71
rect 33 31 2025 37
rect -2025 -37 -33 -31
rect -2025 -71 -2013 -37
rect -45 -71 -33 -37
rect -2025 -77 -33 -71
rect 33 -37 2025 -31
rect 33 -71 45 -37
rect 2013 -71 2025 -37
rect 33 -77 2025 -71
rect -2081 -130 -2035 -118
rect -2081 -2106 -2075 -130
rect -2041 -2106 -2035 -130
rect -2081 -2118 -2035 -2106
rect -23 -130 23 -118
rect -23 -2106 -17 -130
rect 17 -2106 23 -130
rect -23 -2118 23 -2106
rect 2035 -130 2081 -118
rect 2035 -2106 2041 -130
rect 2075 -2106 2081 -130
rect 2035 -2118 2081 -2106
rect -2025 -2165 -33 -2159
rect -2025 -2199 -2013 -2165
rect -45 -2199 -33 -2165
rect -2025 -2205 -33 -2199
rect 33 -2165 2025 -2159
rect 33 -2199 45 -2165
rect 2013 -2199 2025 -2165
rect 33 -2205 2025 -2199
<< properties >>
string FIXED_BBOX -2172 -2284 2172 2284
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 10 l 10.0 m 2 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
