magic
tech sky130A
magscale 1 2
timestamp 1713128983
<< error_s >>
rect 10100 300 10106 306
rect 10094 294 10100 300
rect 10094 100 10100 106
rect 10300 100 10306 106
rect 10100 94 10106 100
rect 10294 94 10300 100
rect 8600 -1000 8606 -994
rect 8794 -1000 8800 -994
rect 8594 -1006 8600 -1000
rect 8800 -1006 8806 -1000
rect 8594 -1200 8600 -1194
rect 8800 -1200 8806 -1194
rect 8600 -1206 8606 -1200
rect 8794 -1206 8800 -1200
rect 7100 -2400 7106 -2394
rect 7294 -2400 7300 -2394
rect 7094 -2406 7100 -2400
rect 7300 -2406 7306 -2400
rect 7094 -2600 7100 -2594
rect 7300 -2600 7306 -2594
rect 7100 -2606 7106 -2600
rect 7294 -2606 7300 -2600
<< locali >>
rect 6500 4494 6900 4500
rect 6500 4306 6606 4494
rect 6794 4306 6900 4494
rect 6500 4300 6900 4306
rect 8200 4495 8700 4500
rect 8200 4305 8305 4495
rect 8495 4305 8700 4495
rect 8200 4300 8700 4305
<< viali >>
rect 6606 4306 6794 4494
rect 8305 4305 8495 4495
<< metal1 >>
rect 7400 4800 7600 4806
rect 5694 4600 5700 4800
rect 5900 4600 5906 4800
rect 7400 4594 7600 4600
rect 6580 4494 6820 4520
rect 6580 4306 6606 4494
rect 6794 4306 6820 4494
rect 6580 4280 6820 4306
rect 8299 4495 8501 4507
rect 9294 4500 9300 4700
rect 9500 4500 9506 4700
rect 10294 4500 10300 4700
rect 10500 4500 10506 4700
rect 8299 4305 8305 4495
rect 8495 4305 8501 4495
rect 5200 3800 5400 3806
rect 6600 3800 6800 4280
rect 7900 3800 8100 3806
rect 6300 3600 7000 3800
rect 5200 3594 5400 3600
rect 6600 2200 6800 3600
rect 7900 3594 8100 3600
rect 8299 2201 8501 4305
rect 10699 2201 10901 2207
rect 8299 2200 8799 2201
rect 5100 2000 8799 2200
rect 8299 1999 8799 2000
rect 9001 1999 9007 2201
rect 10699 1993 10901 1999
rect 5100 1700 7000 1900
rect 5100 1400 6700 1600
rect 5680 300 5920 320
rect 5680 100 5700 300
rect 5900 100 5920 300
rect 5680 80 5920 100
rect 5180 -600 5420 -580
rect 5180 -800 5200 -600
rect 5400 -800 5420 -600
rect 5180 -820 5420 -800
rect 6100 -600 6300 -594
rect 6100 -806 6300 -800
rect 5400 -1200 5600 -900
rect 5900 -1200 6100 -900
rect 6500 -1200 6700 1400
rect 5400 -1400 6700 -1200
rect 6800 -1200 7000 1700
rect 9000 1400 9200 1800
rect 9600 1400 10000 1500
rect 9000 1200 9700 1400
rect 9900 1200 10000 1400
rect 9600 1100 10000 1200
rect 7594 100 7600 300
rect 7800 100 7806 300
rect 10300 100 11100 300
rect 8000 -600 8200 -594
rect 7094 -800 7100 -600
rect 7300 -800 7306 -600
rect 8000 -806 8200 -800
rect 7300 -1200 7500 -900
rect 7800 -1200 8000 -900
rect 8900 -1200 9400 -1000
rect 6800 -1400 8000 -1200
rect 5400 -1700 5600 -1400
rect 5900 -1700 6100 -1400
rect 7300 -1700 7500 -1400
rect 7800 -1700 8000 -1400
rect 8760 -1700 8980 -1640
rect 5600 -2000 5800 -1994
rect 5600 -2206 5800 -2200
rect 7500 -2000 7700 -1994
rect 7500 -2206 7700 -2200
rect 6000 -2400 6200 -2394
rect 7900 -2400 8100 -2394
rect 5194 -2600 5200 -2400
rect 5400 -2600 5406 -2400
rect 8700 -2500 8900 -1700
rect 9100 -1900 9106 -1700
rect 9200 -2300 9400 -1200
rect 10100 -1700 10300 100
rect 9900 -1900 10300 -1700
rect 9000 -2500 9700 -2300
rect 6000 -2606 6200 -2600
rect 7900 -2606 8100 -2600
rect 8300 -2700 8900 -2500
rect 8300 -2900 8500 -2700
rect 9200 -2900 9400 -2500
rect 9700 -2700 9900 -2618
rect 9694 -2897 9700 -2700
rect 9900 -2897 9906 -2700
<< via1 >>
rect 5700 4600 5900 4800
rect 7400 4600 7600 4800
rect 9300 4500 9500 4700
rect 10300 4500 10500 4700
rect 5200 3600 5400 3800
rect 7900 3600 8100 3800
rect 8799 1999 9001 2201
rect 10699 1999 10901 2201
rect 5700 100 5900 300
rect 5200 -800 5400 -600
rect 6100 -800 6300 -600
rect 9700 1200 9900 1400
rect 7600 100 7800 300
rect 10100 100 10300 300
rect 7100 -800 7300 -600
rect 8000 -800 8200 -600
rect 8600 -1200 8800 -1000
rect 5600 -2200 5800 -2000
rect 7500 -2200 7700 -2000
rect 5200 -2600 5400 -2400
rect 6000 -2600 6200 -2400
rect 7100 -2600 7300 -2400
rect 7900 -2600 8100 -2400
rect 8900 -1900 9100 -1700
rect 9700 -2897 9900 -2700
<< metal2 >>
rect 5700 4800 5900 4806
rect 5900 4600 7400 4800
rect 7600 4600 7606 4800
rect 9300 4700 9500 4706
rect 5700 3800 5900 4600
rect 9300 3800 9500 4500
rect 10300 4700 10500 4706
rect 10300 3800 10500 4500
rect 5194 3600 5200 3800
rect 5400 3600 5900 3800
rect 5700 320 5900 3600
rect 7600 3600 7900 3800
rect 8100 3600 10500 3800
rect 5680 300 5920 320
rect 5680 100 5700 300
rect 5900 100 5920 300
rect 5680 80 5920 100
rect 7600 300 7800 3600
rect 8799 2201 9001 2207
rect 9001 1999 10699 2201
rect 10901 1999 10907 2201
rect 8799 1993 9001 1999
rect 9694 1200 9700 1400
rect 9900 1200 10300 1400
rect 10100 300 10300 1200
rect 7600 94 7800 100
rect 5180 -600 5420 -580
rect 7100 -600 7300 -594
rect 5100 -800 5200 -600
rect 5400 -800 6100 -600
rect 6300 -800 6306 -600
rect 7300 -800 8000 -600
rect 5100 -820 5420 -800
rect 7100 -806 7300 -800
rect 5100 -2000 5300 -820
rect 8200 -2000 8400 -600
rect 5100 -2200 5600 -2000
rect 5800 -2200 5806 -2000
rect 7494 -2200 7500 -2000
rect 7700 -2200 8400 -2000
rect 8500 -1200 8600 -1000
rect 5200 -2400 5400 -2394
rect 8500 -2400 8700 -1200
rect 8900 -1700 9100 -1694
rect 9100 -1900 9700 -1700
rect 8900 -1906 9100 -1900
rect 5400 -2600 6000 -2400
rect 6200 -2600 7100 -2400
rect 7300 -2600 7900 -2400
rect 8100 -2600 8700 -2400
rect 5200 -2606 5400 -2600
rect 9500 -2694 9700 -1900
rect 9500 -2700 9900 -2694
rect 9500 -2897 9700 -2700
rect 9500 -2900 9900 -2897
rect 9700 -2903 9900 -2900
use sky130_fd_pr__cap_mim_m3_1_VCAG9S  XC2
timestamp 1713045697
transform -1 0 7686 0 -1 1940
box -686 -540 686 540
use sky130_fd_pr__nfet_01v8_QGMQL3  XM1
timestamp 1713045697
transform 1 0 8872 0 1 -2374
box -296 -460 296 460
use sky130_fd_pr__nfet_01v8_MMMA4V  XM2
timestamp 1713045697
transform 1 0 8872 0 1 -1100
box -296 -710 296 710
use sky130_fd_pr__nfet_01v8_HS3BL4  XM3
timestamp 1713045697
transform 1 0 9796 0 1 -1790
box -296 -1010 296 1010
use sky130_fd_pr__nfet_01v8_W2FWA4  XM4
timestamp 1713050122
transform 1 0 5725 0 1 -2190
box -625 -710 625 710
use sky130_fd_pr__nfet_01v8_J222PV  XM5
timestamp 1713050122
transform 1 0 7625 0 1 -2190
box -625 -710 625 710
use sky130_fd_pr__pfet_01v8_6H4ZLK  XM6
timestamp 1713045697
transform 0 -1 5819 1 0 3696
box -1196 -719 1196 719
use sky130_fd_pr__pfet_01v8_6H4ZLK  XM7
timestamp 1713045697
transform 0 1 7519 -1 0 3696
box -1196 -719 1196 719
use sky130_fd_pr__pfet_01v8_ST5LSM  XM8
timestamp 1713050389
transform 1 0 9825 0 1 2619
box -1225 -2219 1225 2219
use sky130_fd_pr__nfet_05v0_nvt_CXW7PW  XM9
timestamp 1713050122
transform -1 0 5757 0 -1 58
box -657 -1258 657 1258
use sky130_fd_pr__nfet_05v0_nvt_CXW7PW  XM10
timestamp 1713050122
transform 1 0 7657 0 1 58
box -657 -1258 657 1258
<< labels >>
flabel metal1 5100 1400 5300 1600 0 FreeSans 256 0 0 0 vn
port 3 nsew
flabel metal1 5100 1700 5300 1900 0 FreeSans 256 0 0 0 vp
port 2 nsew
flabel metal1 8300 -2900 8500 -2700 0 FreeSans 256 0 0 0 ibias
port 4 nsew
flabel metal1 9200 -2900 9400 -2700 0 FreeSans 256 0 0 0 vss
port 5 nsew
flabel metal1 5100 2000 5300 2200 0 FreeSans 256 0 0 0 vdd
port 0 nsew
flabel metal1 10900 100 11100 300 0 FreeSans 256 0 0 0 vo
port 1 nsew
<< end >>
