magic
tech sky130A
magscale 1 2
timestamp 1713051387
<< pwell >>
rect -1054 -927 1054 927
<< psubdiff >>
rect -1018 857 -922 891
rect 922 857 1018 891
rect -1018 795 -984 857
rect 984 795 1018 857
rect -1018 -857 -984 -795
rect 984 -857 1018 -795
rect -1018 -891 -922 -857
rect 922 -891 1018 -857
<< psubdiffcont >>
rect -922 857 922 891
rect -1018 -795 -984 795
rect 984 -795 1018 795
rect -922 -891 922 -857
<< xpolycontact >>
rect -888 329 -750 761
rect -888 -761 -750 -329
rect -654 329 -516 761
rect -654 -761 -516 -329
rect -420 329 -282 761
rect -420 -761 -282 -329
rect -186 329 -48 761
rect -186 -761 -48 -329
rect 48 329 186 761
rect 48 -761 186 -329
rect 282 329 420 761
rect 282 -761 420 -329
rect 516 329 654 761
rect 516 -761 654 -329
rect 750 329 888 761
rect 750 -761 888 -329
<< xpolyres >>
rect -888 -329 -750 329
rect -654 -329 -516 329
rect -420 -329 -282 329
rect -186 -329 -48 329
rect 48 -329 186 329
rect 282 -329 420 329
rect 516 -329 654 329
rect 750 -329 888 329
<< locali >>
rect -1018 857 -922 891
rect 922 857 1018 891
rect -1018 795 -984 857
rect 984 795 1018 857
rect -1018 -857 -984 -795
rect 984 -857 1018 -795
rect -1018 -891 -922 -857
rect 922 -891 1018 -857
<< viali >>
rect -872 346 -766 743
rect -638 346 -532 743
rect -404 346 -298 743
rect -170 346 -64 743
rect 64 346 170 743
rect 298 346 404 743
rect 532 346 638 743
rect 766 346 872 743
rect -872 -743 -766 -346
rect -638 -743 -532 -346
rect -404 -743 -298 -346
rect -170 -743 -64 -346
rect 64 -743 170 -346
rect 298 -743 404 -346
rect 532 -743 638 -346
rect 766 -743 872 -346
<< metal1 >>
rect -878 743 -760 755
rect -878 346 -872 743
rect -766 346 -760 743
rect -878 334 -760 346
rect -644 743 -526 755
rect -644 346 -638 743
rect -532 346 -526 743
rect -644 334 -526 346
rect -410 743 -292 755
rect -410 346 -404 743
rect -298 346 -292 743
rect -410 334 -292 346
rect -176 743 -58 755
rect -176 346 -170 743
rect -64 346 -58 743
rect -176 334 -58 346
rect 58 743 176 755
rect 58 346 64 743
rect 170 346 176 743
rect 58 334 176 346
rect 292 743 410 755
rect 292 346 298 743
rect 404 346 410 743
rect 292 334 410 346
rect 526 743 644 755
rect 526 346 532 743
rect 638 346 644 743
rect 526 334 644 346
rect 760 743 878 755
rect 760 346 766 743
rect 872 346 878 743
rect 760 334 878 346
rect -878 -346 -760 -334
rect -878 -743 -872 -346
rect -766 -743 -760 -346
rect -878 -755 -760 -743
rect -644 -346 -526 -334
rect -644 -743 -638 -346
rect -532 -743 -526 -346
rect -644 -755 -526 -743
rect -410 -346 -292 -334
rect -410 -743 -404 -346
rect -298 -743 -292 -346
rect -410 -755 -292 -743
rect -176 -346 -58 -334
rect -176 -743 -170 -346
rect -64 -743 -58 -346
rect -176 -755 -58 -743
rect 58 -346 176 -334
rect 58 -743 64 -346
rect 170 -743 176 -346
rect 58 -755 176 -743
rect 292 -346 410 -334
rect 292 -743 298 -346
rect 404 -743 410 -346
rect 292 -755 410 -743
rect 526 -346 644 -334
rect 526 -743 532 -346
rect 638 -743 644 -346
rect 526 -755 644 -743
rect 760 -346 878 -334
rect 760 -743 766 -346
rect 872 -743 878 -346
rect 760 -755 878 -743
<< properties >>
string FIXED_BBOX -1001 -874 1001 874
string gencell sky130_fd_pr__res_xhigh_po_0p69
string library sky130
string parameters w 0.690 l 3.45 m 1 nx 8 wmin 0.690 lmin 0.50 rho 2000 val 10.545k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.690 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
