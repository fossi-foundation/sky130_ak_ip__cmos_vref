magic
tech sky130A
magscale 1 2
timestamp 1717344711
<< metal1 >>
rect 700 -300 2894 -100
rect 2044 -558 2436 -300
rect 2502 -558 2894 -300
rect 835 -602 899 -590
rect 835 -1578 841 -602
rect 893 -1578 899 -602
rect 835 -1590 899 -1578
rect 1040 -1622 1140 -558
rect 1292 -960 1356 -590
rect 1200 -980 1440 -960
rect 1200 -1180 1220 -980
rect 1420 -1180 1440 -980
rect 1200 -1200 1440 -1180
rect 1292 -1590 1356 -1200
rect 1500 -1622 1600 -558
rect 1751 -602 1815 -590
rect 1751 -866 1757 -602
rect 1809 -866 1815 -602
rect 1751 -1316 1815 -866
rect 1751 -1580 1757 -1316
rect 1809 -1580 1815 -1316
rect 1751 -1590 1815 -1580
rect 1979 -1316 2043 -590
rect 1979 -1580 1985 -1316
rect 2037 -1580 2043 -1316
rect 1979 -1590 2043 -1580
rect 900 -1800 1292 -1622
rect 1358 -1800 1750 -1622
rect 2180 -1640 2280 -558
rect 2437 -960 2501 -590
rect 2360 -980 2600 -960
rect 2360 -1180 2380 -980
rect 2580 -1180 2600 -980
rect 2360 -1200 2600 -1180
rect 2437 -1594 2501 -1200
rect 2680 -1640 2780 -558
rect 2894 -604 2958 -590
rect 2894 -866 2900 -604
rect 2952 -866 2958 -604
rect 2894 -1308 2958 -866
rect 2894 -1580 2900 -1308
rect 2952 -1580 2958 -1308
rect 2894 -1590 2958 -1580
rect 700 -2000 1750 -1800
rect 700 -2300 1750 -2100
rect 900 -2458 1292 -2300
rect 1358 -2458 1750 -2300
rect 3100 -2180 3300 -100
rect 3560 -300 3800 -100
rect 3560 -320 3720 -300
rect 3560 -720 3580 -320
rect 3700 -720 3720 -320
rect 3560 -760 3720 -720
rect 3920 -760 4320 -300
rect 4520 -760 4920 -300
rect 4980 -760 5380 -300
rect 3560 -1420 4080 -1400
rect 3560 -1820 3580 -1420
rect 3700 -1820 4080 -1420
rect 3560 -1840 4080 -1820
rect 4160 -1420 4680 -1400
rect 4160 -1820 4180 -1420
rect 4300 -1820 4680 -1420
rect 4160 -1840 4680 -1820
rect 4760 -1840 5140 -1400
rect 5220 -1420 5380 -1400
rect 5220 -1820 5240 -1420
rect 5360 -1820 5380 -1420
rect 5220 -1840 5380 -1820
rect 3100 -2420 3720 -2180
rect 834 -2504 898 -2490
rect 834 -2766 840 -2504
rect 892 -2766 898 -2504
rect 834 -3216 898 -2766
rect 834 -3480 840 -3216
rect 892 -3480 898 -3216
rect 834 -3490 898 -3480
rect 1040 -3540 1140 -2458
rect 1293 -2880 1357 -2490
rect 1200 -2900 1440 -2880
rect 1200 -3100 1220 -2900
rect 1420 -3100 1440 -2900
rect 1200 -3120 1440 -3100
rect 1293 -3490 1357 -3120
rect 1500 -3540 1600 -2458
rect 1751 -2504 1815 -2490
rect 1751 -2766 1757 -2504
rect 1809 -2766 1815 -2504
rect 1751 -3216 1815 -2766
rect 1751 -3480 1757 -3216
rect 1809 -3480 1815 -3216
rect 1751 -3490 1815 -3480
rect 1979 -2504 2043 -2488
rect 1979 -2766 1985 -2504
rect 2037 -2766 2043 -2504
rect 1979 -3216 2043 -2766
rect 1979 -3480 1985 -3216
rect 2037 -3480 2043 -3216
rect 1979 -3490 2043 -3480
rect 2200 -3522 2300 -2440
rect 2438 -2880 2502 -2490
rect 2360 -2900 2600 -2880
rect 2360 -3100 2380 -2900
rect 2580 -3100 2600 -2900
rect 2360 -3120 2600 -3100
rect 2438 -3490 2502 -3120
rect 2660 -3522 2760 -2440
rect 2896 -2504 2960 -2490
rect 2896 -2766 2902 -2504
rect 2954 -2766 2960 -2504
rect 3300 -2620 3720 -2420
rect 3100 -2640 3720 -2620
rect 3780 -2640 4180 -2180
rect 4260 -2640 4660 -2180
rect 4720 -2640 5120 -2180
rect 5200 -2200 5360 -2180
rect 5200 -2620 5220 -2200
rect 5340 -2620 5360 -2200
rect 5200 -2640 5360 -2620
rect 2896 -3216 2960 -2766
rect 2896 -3480 2902 -3216
rect 2954 -3480 2960 -3216
rect 2896 -3490 2960 -3480
rect 2044 -3700 2436 -3522
rect 2502 -3700 2894 -3522
rect 700 -3900 2894 -3700
rect 3560 -3720 3940 -3280
rect 4020 -3720 4420 -3280
rect 4500 -3720 4880 -3280
rect 4960 -3720 5360 -3280
<< via1 >>
rect 841 -1578 893 -602
rect 1220 -1180 1420 -980
rect 1757 -866 1809 -602
rect 1757 -1580 1809 -1316
rect 1985 -1580 2037 -1316
rect 2380 -1180 2580 -980
rect 2900 -866 2952 -604
rect 2900 -1580 2952 -1308
rect 3580 -720 3700 -320
rect 3580 -1820 3700 -1420
rect 4180 -1820 4300 -1420
rect 5240 -1820 5360 -1420
rect 840 -2766 892 -2504
rect 840 -3480 892 -3216
rect 1220 -3100 1420 -2900
rect 1757 -2766 1809 -2504
rect 1757 -3480 1809 -3216
rect 1985 -2766 2037 -2504
rect 1985 -3480 2037 -3216
rect 2380 -3100 2580 -2900
rect 2902 -2766 2954 -2504
rect 3100 -2620 3300 -2420
rect 5220 -2620 5340 -2200
rect 2902 -3480 2954 -3216
<< metal2 >>
rect 3560 -320 3720 -300
rect 835 -602 899 -590
rect 835 -1578 841 -602
rect 893 -640 899 -602
rect 1751 -602 1815 -590
rect 1751 -640 1757 -602
rect 893 -840 1757 -640
rect 893 -1340 899 -840
rect 1751 -866 1757 -840
rect 1809 -640 1815 -602
rect 2894 -604 2958 -590
rect 1809 -840 2580 -640
rect 1809 -866 1815 -840
rect 1751 -872 1815 -866
rect 2380 -960 2580 -840
rect 2894 -866 2900 -604
rect 2952 -640 2958 -604
rect 3560 -640 3580 -320
rect 2952 -720 3580 -640
rect 3700 -720 3720 -320
rect 2952 -840 3720 -720
rect 2952 -866 2958 -840
rect 2894 -877 2958 -866
rect 1200 -980 1440 -960
rect 2360 -980 2600 -960
rect 1200 -1180 1220 -980
rect 1420 -1180 1945 -980
rect 1200 -1200 1440 -1180
rect 1751 -1316 1815 -1308
rect 1751 -1340 1757 -1316
rect 893 -1540 1757 -1340
rect 893 -1578 899 -1540
rect 835 -1590 899 -1578
rect 1751 -1580 1757 -1540
rect 1809 -1580 1815 -1316
rect 1751 -1590 1815 -1580
rect 1845 -1800 1945 -1180
rect 2360 -1180 2380 -980
rect 2580 -1180 3720 -980
rect 2360 -1200 2600 -1180
rect 2894 -1308 2958 -1300
rect 1979 -1316 2043 -1308
rect 1979 -1580 1985 -1316
rect 2037 -1340 2043 -1316
rect 2894 -1340 2900 -1308
rect 2037 -1540 2900 -1340
rect 2037 -1580 2043 -1540
rect 1979 -1590 2043 -1580
rect 2894 -1580 2900 -1540
rect 2952 -1580 2958 -1308
rect 2894 -1590 2958 -1580
rect 3560 -1420 3720 -1180
rect 1845 -1880 3520 -1800
rect 3560 -1820 3580 -1420
rect 3700 -1820 3720 -1420
rect 3560 -1840 3720 -1820
rect 4160 -1420 4320 -1400
rect 4160 -1820 4180 -1420
rect 4300 -1820 4320 -1420
rect 4160 -1880 4320 -1820
rect 1845 -2000 4320 -1880
rect 5220 -1420 5380 -1400
rect 5220 -1820 5240 -1420
rect 5360 -1820 5380 -1420
rect 1845 -2490 1945 -2000
rect 5220 -2040 5380 -1820
rect 2820 -2180 5380 -2040
rect 834 -2504 898 -2490
rect 834 -2766 840 -2504
rect 892 -2540 898 -2504
rect 1751 -2504 1945 -2490
rect 1751 -2540 1757 -2504
rect 892 -2740 1757 -2540
rect 892 -2766 898 -2740
rect 834 -3216 898 -2766
rect 1751 -2766 1757 -2740
rect 1809 -2766 1945 -2504
rect 1751 -2778 1945 -2766
rect 1979 -2504 2043 -2488
rect 1979 -2766 1985 -2504
rect 2037 -2520 2043 -2504
rect 2820 -2504 2960 -2180
rect 5200 -2200 5360 -2180
rect 2820 -2520 2902 -2504
rect 2037 -2720 2902 -2520
rect 2037 -2766 2043 -2720
rect 1200 -2900 1440 -2880
rect 1979 -2900 2043 -2766
rect 2896 -2766 2902 -2720
rect 2954 -2766 2960 -2504
rect 2896 -2778 2960 -2766
rect 3100 -2420 3300 -2414
rect 1200 -3100 1220 -2900
rect 1420 -3100 2043 -2900
rect 1200 -3120 1440 -3100
rect 834 -3480 840 -3216
rect 892 -3240 898 -3216
rect 1751 -3216 1815 -3202
rect 1751 -3240 1757 -3216
rect 892 -3440 1757 -3240
rect 892 -3480 898 -3440
rect 834 -3490 898 -3480
rect 1751 -3480 1757 -3440
rect 1809 -3480 1815 -3216
rect 1751 -3490 1815 -3480
rect 1979 -3216 2043 -3100
rect 2360 -2900 2600 -2880
rect 3100 -2900 3300 -2620
rect 5200 -2620 5220 -2200
rect 5340 -2620 5360 -2200
rect 5200 -2640 5360 -2620
rect 2360 -3100 2380 -2900
rect 2580 -3100 3300 -2900
rect 2360 -3120 2600 -3100
rect 1979 -3480 1985 -3216
rect 2037 -3240 2043 -3216
rect 2896 -3216 2960 -3202
rect 2896 -3240 2902 -3216
rect 2037 -3440 2902 -3240
rect 2037 -3480 2043 -3440
rect 1979 -3490 2043 -3480
rect 2896 -3480 2902 -3440
rect 2954 -3480 2960 -3216
rect 2896 -3490 2960 -3480
use sky130_fd_pr__res_xhigh_po_0p69_2G52HS  sky130_fd_pr__res_xhigh_po_0p69_2G52HS_0 paramcells
timestamp 1713051387
transform 1 0 4116 0 1 -1073
box -352 -927 352 927
use sky130_fd_pr__res_xhigh_po_0p69_D5BT6X  sky130_fd_pr__res_xhigh_po_0p69_D5BT6X_0 paramcells
timestamp 1713051387
transform 1 0 4454 0 1 -2953
box -1054 -927 1054 927
use sky130_fd_pr__res_xhigh_po_0p69_H5FMR6  sky130_fd_pr__res_xhigh_po_0p69_H5FMR6_0 paramcells
timestamp 1713051387
transform 1 0 3635 0 1 -1073
box -235 -927 235 927
use sky130_fd_pr__res_xhigh_po_0p69_H5TM75  sky130_fd_pr__res_xhigh_po_0p69_H5TM75_0 paramcells
timestamp 1713051387
transform 1 0 4948 0 1 -1073
box -586 -927 586 927
use sky130_fd_pr__nfet_01v8_J222PV  XM1 paramcells
timestamp 1713050122
transform 1 0 2469 0 1 -1090
box -625 -710 625 710
use sky130_fd_pr__nfet_01v8_J222PV  XM2
timestamp 1713050122
transform 1 0 1325 0 1 -1090
box -625 -710 625 710
use sky130_fd_pr__nfet_01v8_J222PV  XM3
timestamp 1713050122
transform 1 0 1325 0 1 -2990
box -625 -710 625 710
use sky130_fd_pr__nfet_01v8_J222PV  XM4
timestamp 1713050122
transform 1 0 2469 0 1 -2990
box -625 -710 625 710
<< labels >>
flabel metal1 700 -2000 900 -1800 0 FreeSans 256 0 0 0 trim1
port 5 nsew
flabel metal1 700 -2300 900 -2100 0 FreeSans 256 0 0 0 trim2
port 3 nsew
flabel metal1 700 -3900 900 -3700 0 FreeSans 256 0 0 0 trim3
port 4 nsew
flabel metal1 3100 -300 3300 -100 0 FreeSans 256 0 0 0 A
port 1 nsew
flabel metal1 700 -300 900 -100 0 FreeSans 256 0 0 0 trim0
port 2 nsew
flabel metal1 3600 -300 3800 -100 0 FreeSans 256 0 0 0 B
port 6 nsew
<< end >>
