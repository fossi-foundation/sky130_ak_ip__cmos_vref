magic
tech sky130A
magscale 1 2
timestamp 1716339083
<< dnwell >>
rect 8800 -19700 21700 0
<< nwell >>
rect 8720 -1800 21780 80
rect 8720 -19494 9006 -1800
rect 21494 -15000 21780 -1800
rect 19000 -17100 21780 -15000
rect 15500 -19494 21780 -17100
rect 8720 -19780 21780 -19494
<< psubdiff >>
rect 21100 -9500 21300 -9476
rect 21100 -9724 21300 -9700
<< nsubdiff >>
rect 8757 23 21743 43
rect 8757 -11 8837 23
rect 21663 -11 21743 23
rect 8757 -31 21743 -11
rect 8757 -37 8831 -31
rect 8757 -19663 8777 -37
rect 8811 -19663 8831 -37
rect 21669 -37 21743 -31
rect 8757 -19669 8831 -19663
rect 21669 -19663 21689 -37
rect 21723 -19663 21743 -37
rect 21669 -19669 21743 -19663
rect 8757 -19689 21743 -19669
rect 8757 -19723 8837 -19689
rect 21663 -19723 21743 -19689
rect 8757 -19743 21743 -19723
<< psubdiffcont >>
rect 21100 -9700 21300 -9500
<< nsubdiffcont >>
rect 8837 -11 21663 23
rect 8777 -19663 8811 -37
rect 21689 -19663 21723 -37
rect 8837 -19723 21663 -19689
<< locali >>
rect 8777 -11 8837 23
rect 21663 -11 21723 23
rect 8777 -37 8811 -11
rect 21689 -37 21723 -11
rect 10953 -8427 10987 -8393
rect 21100 -9500 21300 -9484
rect 21100 -9716 21300 -9700
rect 8777 -19689 8811 -19663
rect 21689 -19689 21723 -19663
rect 8777 -19723 8837 -19689
rect 21663 -19723 21723 -19689
<< viali >>
rect 9667 -8631 9701 -8597
rect 9943 -8631 9977 -8597
rect 10219 -8631 10253 -8597
rect 10495 -8631 10529 -8597
rect 10771 -8631 10805 -8597
rect 9849 -8767 9883 -8733
rect 10125 -8767 10159 -8733
rect 10401 -8767 10435 -8733
rect 10677 -8767 10711 -8733
rect 10953 -8767 10987 -8733
rect 9432 -9932 13966 -9898
rect 9336 -10668 9370 -9994
rect 9336 -11868 9370 -10960
rect 9336 -15368 9370 -12120
<< metal1 >>
rect 8720 -120 21780 80
rect 8720 -6100 8920 -120
rect 9219 -400 14900 -200
rect 9068 -4238 9132 -450
rect 9219 -2449 11719 -2443
rect 9219 -2501 9225 -2449
rect 11713 -2501 11719 -2449
rect 9219 -2507 11719 -2501
rect 9068 -4482 9074 -4238
rect 9126 -4482 9132 -4238
rect 9068 -4488 9132 -4482
rect 11805 -4250 11869 -450
rect 11955 -2449 14455 -2443
rect 11955 -2501 11961 -2449
rect 14449 -2501 14455 -2449
rect 11955 -2507 14455 -2501
rect 11805 -4494 11811 -4250
rect 11863 -4494 11869 -4250
rect 14542 -4238 14606 -450
rect 14542 -4482 14548 -4238
rect 14600 -4482 14606 -4238
rect 14542 -4488 14606 -4482
rect 14700 -3400 14900 -400
rect 15500 -1700 16000 -1500
rect 15500 -3400 15700 -1700
rect 14700 -3600 15700 -3400
rect 11805 -4500 11869 -4494
rect 9219 -4620 11719 -4556
rect 11955 -4620 14455 -4556
rect 14700 -4620 14900 -3600
rect 15000 -3700 15200 -3694
rect 15200 -3900 15400 -3700
rect 15000 -3906 15400 -3900
rect 15200 -4280 15400 -3906
rect 15180 -4300 15420 -4280
rect 15180 -4500 15200 -4300
rect 15400 -4500 15420 -4300
rect 15180 -4520 15420 -4500
rect 9220 -4820 14900 -4620
rect 14877 -4899 15117 -4878
rect 14877 -4900 14900 -4899
rect 9300 -5012 14900 -4900
rect 8999 -5590 9290 -5089
rect 13348 -5400 13412 -5090
rect 14877 -5099 14900 -5012
rect 15100 -4900 15117 -4899
rect 15200 -4900 15400 -4520
rect 15100 -5099 15400 -4900
rect 14877 -5100 15400 -5099
rect 14877 -5122 15117 -5100
rect 15180 -5400 15420 -5380
rect 13348 -5590 15200 -5400
rect 9000 -5800 9200 -5590
rect 13400 -5600 15200 -5590
rect 15400 -5600 15420 -5400
rect 14210 -5652 14410 -5600
rect 15180 -5620 15420 -5600
rect 9300 -5732 14178 -5668
rect 9000 -6000 12100 -5800
rect 12300 -6000 12306 -5800
rect 11945 -6091 13619 -6088
rect 8720 -6300 11619 -6100
rect 11800 -6152 13619 -6091
rect 11800 -6158 12689 -6152
rect 9000 -6600 9200 -6300
rect 9522 -6348 9588 -6341
rect 9522 -6400 9529 -6348
rect 9581 -6400 9588 -6348
rect 9522 -6407 9588 -6400
rect 11650 -6347 11716 -6341
rect 11650 -6399 11657 -6347
rect 11709 -6399 11716 -6347
rect 11650 -6407 11716 -6399
rect 9619 -6500 11619 -6456
rect 11800 -6500 12000 -6158
rect 9619 -6700 12000 -6500
rect 9000 -7040 9200 -6900
rect 10756 -7040 10820 -7038
rect 9000 -7044 10820 -7040
rect 9000 -7096 10762 -7044
rect 10814 -7096 10820 -7044
rect 9000 -7100 10820 -7096
rect 10756 -7102 10820 -7100
rect 9000 -7340 9200 -7200
rect 10480 -7340 10544 -7338
rect 9000 -7344 10544 -7340
rect 9000 -7396 10486 -7344
rect 10538 -7396 10544 -7344
rect 9000 -7400 10544 -7396
rect 10480 -7402 10544 -7400
rect 9000 -7640 9200 -7500
rect 10204 -7640 10268 -7638
rect 9000 -7644 10268 -7640
rect 9000 -7696 10210 -7644
rect 10262 -7696 10268 -7644
rect 9000 -7700 10268 -7696
rect 10204 -7702 10268 -7700
rect 9000 -7940 9200 -7800
rect 9929 -7940 9993 -7938
rect 9000 -7944 9993 -7940
rect 9000 -7996 9935 -7944
rect 9987 -7996 9993 -7944
rect 9000 -8000 9993 -7996
rect 9929 -8002 9993 -8000
rect 9652 -8100 9716 -8098
rect 9000 -8104 9716 -8100
rect 9000 -8156 9658 -8104
rect 9710 -8156 9716 -8104
rect 9000 -8160 9716 -8156
rect 9000 -8300 9200 -8160
rect 9652 -8162 9716 -8160
rect 9500 -8356 9638 -8260
rect 9500 -8400 9596 -8356
rect 9000 -8496 9596 -8400
rect 10938 -8390 11002 -8384
rect 10938 -8442 10944 -8390
rect 10996 -8442 11002 -8390
rect 10938 -8448 11002 -8442
rect 9000 -8600 9200 -8496
rect 9652 -8588 9716 -8582
rect 9652 -8640 9658 -8588
rect 9710 -8640 9716 -8588
rect 9652 -8646 9716 -8640
rect 9929 -8589 9993 -8583
rect 9929 -8641 9935 -8589
rect 9987 -8641 9993 -8589
rect 9929 -8647 9993 -8641
rect 10204 -8588 10268 -8582
rect 10204 -8640 10210 -8588
rect 10262 -8640 10268 -8588
rect 10204 -8646 10268 -8640
rect 10480 -8588 10544 -8582
rect 10480 -8640 10486 -8588
rect 10538 -8640 10544 -8588
rect 10480 -8646 10544 -8640
rect 10756 -8588 10820 -8582
rect 10756 -8640 10762 -8588
rect 10814 -8640 10820 -8588
rect 10756 -8646 10820 -8640
rect 11800 -8600 12000 -6700
rect 12468 -6214 12532 -6208
rect 12468 -8194 12474 -6214
rect 12526 -8194 12532 -6214
rect 12468 -8200 12532 -8194
rect 13706 -6214 13770 -6208
rect 13706 -8194 13712 -6214
rect 13764 -8194 13770 -6214
rect 14068 -7756 14132 -5732
rect 14488 -7756 14552 -5708
rect 14068 -7800 14552 -7756
rect 14068 -8000 14900 -7800
rect 15100 -8000 15106 -7800
rect 13706 -8200 13770 -8194
rect 12619 -8300 13619 -8256
rect 15180 -8300 15420 -8280
rect 12619 -8352 15200 -8300
rect 12700 -8500 15200 -8352
rect 15400 -8500 15420 -8300
rect 15180 -8520 15420 -8500
rect 14580 -8600 14820 -8580
rect 15500 -8600 15700 -3600
rect 15800 -4000 16000 -1800
rect 15800 -4206 16000 -4200
rect 15800 -4300 16000 -4294
rect 15800 -4506 16000 -4500
rect 15780 -5400 16020 -5380
rect 15780 -5600 15800 -5400
rect 16000 -5600 16020 -5400
rect 15780 -5620 16020 -5600
rect 9000 -8804 9200 -8700
rect 9835 -8718 9899 -8712
rect 9835 -8770 9841 -8718
rect 9893 -8770 9899 -8718
rect 9835 -8776 9899 -8770
rect 10111 -8718 10175 -8712
rect 10111 -8770 10117 -8718
rect 10169 -8770 10175 -8718
rect 10111 -8776 10175 -8770
rect 10387 -8718 10451 -8712
rect 10387 -8770 10393 -8718
rect 10445 -8770 10451 -8718
rect 10387 -8776 10451 -8770
rect 10663 -8718 10727 -8712
rect 10663 -8770 10669 -8718
rect 10721 -8770 10727 -8718
rect 10663 -8776 10727 -8770
rect 10939 -8733 11003 -8712
rect 10939 -8767 10953 -8733
rect 10987 -8767 11003 -8733
rect 10939 -8776 11003 -8767
rect 11800 -8800 14600 -8600
rect 14800 -8800 15700 -8600
rect 15800 -8700 16000 -5620
rect 9000 -8900 9638 -8804
rect 14580 -8820 14820 -8800
rect 15800 -8900 19000 -8700
rect 19200 -8900 19206 -8700
rect 10118 -8946 10182 -8940
rect 10118 -8980 10124 -8946
rect 9060 -8998 10124 -8980
rect 10176 -8998 10182 -8946
rect 9060 -9004 10182 -8998
rect 9060 -9040 10180 -9004
rect 8720 -19580 8920 -9100
rect 9060 -17772 9120 -9040
rect 10670 -9100 10730 -9094
rect 9180 -9160 10670 -9100
rect 9180 -15770 9240 -9160
rect 10670 -9166 10730 -9160
rect 14280 -9500 14520 -9480
rect 19600 -9482 19800 -8679
rect 21580 -9101 21780 -120
rect 21094 -9301 21100 -9101
rect 21300 -9301 21780 -9101
rect 19578 -9500 19816 -9482
rect 12080 -9700 12100 -9500
rect 12300 -9700 14300 -9500
rect 14500 -9700 19600 -9500
rect 19800 -9700 21500 -9500
rect 12080 -9862 14100 -9700
rect 14280 -9720 14520 -9700
rect 19578 -9721 19816 -9700
rect 9300 -9880 14100 -9862
rect 9300 -9898 14098 -9880
rect 9300 -9932 9432 -9898
rect 13966 -9932 14098 -9898
rect 9300 -9938 14098 -9932
rect 9300 -9994 9376 -9938
rect 9300 -10668 9336 -9994
rect 9370 -10668 9376 -9994
rect 15194 -10000 15200 -9800
rect 15400 -10000 18700 -9800
rect 18900 -10000 18906 -9800
rect 18994 -10000 19000 -9800
rect 19200 -10000 21500 -9800
rect 9471 -10158 13299 -10040
rect 13925 -10100 14300 -10040
rect 13925 -10158 20500 -10100
rect 13199 -10274 13299 -10158
rect 9471 -10626 9892 -10274
rect 13199 -10392 13925 -10274
rect 14100 -10300 20500 -10158
rect 20700 -10300 21500 -10100
rect 17880 -10400 18120 -10380
rect 14100 -10508 17900 -10400
rect 13925 -10600 17900 -10508
rect 18100 -10600 21500 -10400
rect 13925 -10626 14300 -10600
rect 17880 -10620 18120 -10600
rect 9300 -10960 9376 -10668
rect 9300 -11868 9336 -10960
rect 9370 -11868 9376 -10960
rect 14100 -10900 21500 -10700
rect 14100 -11004 14220 -10900
rect 9472 -11356 9893 -11004
rect 13597 -11122 14220 -11004
rect 15800 -11400 16000 -10900
rect 18700 -11300 19100 -11200
rect 9472 -11824 9893 -11472
rect 17894 -11500 17900 -11300
rect 18100 -11500 18106 -11300
rect 18700 -11500 18800 -11300
rect 19000 -11500 19100 -11300
rect 18700 -11600 19100 -11500
rect 19500 -11300 19900 -11200
rect 19500 -11500 19600 -11300
rect 19800 -11500 19900 -11300
rect 19500 -11600 19900 -11500
rect 20400 -11300 20800 -11200
rect 21094 -11300 21100 -11100
rect 21300 -11300 21800 -11100
rect 20400 -11500 20500 -11300
rect 20700 -11500 20800 -11300
rect 20400 -11600 20800 -11500
rect 14018 -11824 14220 -11706
rect 9300 -12120 9376 -11868
rect 9300 -15368 9336 -12120
rect 9370 -15368 9376 -12120
rect 14100 -12164 14220 -11824
rect 18800 -11908 19000 -11600
rect 19600 -11908 19800 -11600
rect 20500 -11908 20700 -11600
rect 9472 -12516 9893 -12164
rect 13651 -12282 14000 -12164
rect 14072 -12282 15400 -12164
rect 9472 -12984 9893 -12632
rect 13651 -12750 14072 -12398
rect 9472 -13452 9893 -13100
rect 13651 -13218 14072 -12866
rect 14294 -12900 14300 -12700
rect 14500 -12900 14506 -12700
rect 14594 -12900 14600 -12700
rect 14800 -12900 14806 -12700
rect 14894 -12900 14900 -12700
rect 15100 -12900 15106 -12700
rect 9472 -13920 9893 -13568
rect 13651 -13686 14072 -13334
rect 9472 -14388 9893 -14036
rect 13651 -14154 14072 -13802
rect 9472 -14856 9893 -14504
rect 13651 -14622 14072 -14270
rect 9472 -15324 9893 -14972
rect 13651 -15090 14072 -14738
rect 11700 -15324 13772 -15206
rect 9300 -15500 9376 -15368
rect 11700 -15700 11900 -15324
rect 14300 -15500 14500 -12900
rect 12200 -15700 14500 -15500
rect 9180 -15830 9310 -15770
rect 14600 -16608 14800 -12900
rect 14900 -16308 15100 -12900
rect 15200 -16008 15400 -12282
rect 15200 -16208 15700 -16008
rect 14900 -16508 15700 -16308
rect 14600 -16808 15700 -16608
rect 9280 -17400 9520 -17380
rect 9280 -17600 9300 -17400
rect 9500 -17600 9520 -17400
rect 9280 -17620 9520 -17600
rect 9060 -17832 9300 -17772
rect 9280 -19300 9520 -19280
rect 9280 -19500 9300 -19300
rect 9500 -19500 9520 -19300
rect 9280 -19520 9520 -19500
rect 21580 -19580 21780 -11300
rect 8720 -19780 21780 -19580
<< via1 >>
rect 9225 -2501 11713 -2449
rect 9074 -4482 9126 -4238
rect 11961 -2501 14449 -2449
rect 11811 -4494 11863 -4250
rect 14548 -4482 14600 -4238
rect 15000 -3900 15200 -3700
rect 15200 -4500 15400 -4300
rect 14900 -5099 15100 -4899
rect 15200 -5600 15400 -5400
rect 12100 -6000 12300 -5800
rect 9529 -6400 9581 -6348
rect 11657 -6399 11709 -6347
rect 10762 -7096 10814 -7044
rect 10486 -7396 10538 -7344
rect 10210 -7696 10262 -7644
rect 9935 -7996 9987 -7944
rect 9658 -8156 9710 -8104
rect 10944 -8442 10996 -8390
rect 9658 -8597 9710 -8588
rect 9658 -8631 9667 -8597
rect 9667 -8631 9701 -8597
rect 9701 -8631 9710 -8597
rect 9658 -8640 9710 -8631
rect 9935 -8597 9987 -8589
rect 9935 -8631 9943 -8597
rect 9943 -8631 9977 -8597
rect 9977 -8631 9987 -8597
rect 9935 -8641 9987 -8631
rect 10210 -8597 10262 -8588
rect 10210 -8631 10219 -8597
rect 10219 -8631 10253 -8597
rect 10253 -8631 10262 -8597
rect 10210 -8640 10262 -8631
rect 10486 -8597 10538 -8588
rect 10486 -8631 10495 -8597
rect 10495 -8631 10529 -8597
rect 10529 -8631 10538 -8597
rect 10486 -8640 10538 -8631
rect 10762 -8597 10814 -8588
rect 10762 -8631 10771 -8597
rect 10771 -8631 10805 -8597
rect 10805 -8631 10814 -8597
rect 10762 -8640 10814 -8631
rect 12474 -8194 12526 -6214
rect 13712 -8194 13764 -6214
rect 14900 -8000 15100 -7800
rect 15200 -8500 15400 -8300
rect 15800 -4200 16000 -4000
rect 15800 -4500 16000 -4300
rect 15800 -5600 16000 -5400
rect 9841 -8733 9893 -8718
rect 9841 -8767 9849 -8733
rect 9849 -8767 9883 -8733
rect 9883 -8767 9893 -8733
rect 9841 -8770 9893 -8767
rect 10117 -8733 10169 -8718
rect 10117 -8767 10125 -8733
rect 10125 -8767 10159 -8733
rect 10159 -8767 10169 -8733
rect 10117 -8770 10169 -8767
rect 10393 -8733 10445 -8718
rect 10393 -8767 10401 -8733
rect 10401 -8767 10435 -8733
rect 10435 -8767 10445 -8733
rect 10393 -8770 10445 -8767
rect 10669 -8733 10721 -8718
rect 10669 -8767 10677 -8733
rect 10677 -8767 10711 -8733
rect 10711 -8767 10721 -8733
rect 10669 -8770 10721 -8767
rect 14600 -8800 14800 -8600
rect 19000 -8900 19200 -8700
rect 10124 -8998 10176 -8946
rect 10670 -9160 10730 -9100
rect 21100 -9301 21300 -9101
rect 12100 -9700 12300 -9500
rect 14300 -9700 14500 -9500
rect 19600 -9700 19800 -9500
rect 15200 -10000 15400 -9800
rect 18700 -10000 18900 -9800
rect 19000 -10000 19200 -9800
rect 20500 -10300 20700 -10100
rect 17900 -10600 18100 -10400
rect 17900 -11500 18100 -11300
rect 18800 -11500 19000 -11300
rect 19600 -11500 19800 -11300
rect 21100 -11300 21300 -11100
rect 20500 -11500 20700 -11300
rect 14300 -12900 14500 -12700
rect 14600 -12900 14800 -12700
rect 14900 -12900 15100 -12700
rect 9300 -17600 9500 -17400
rect 9300 -19500 9500 -19300
<< metal2 >>
rect 9219 -2449 15200 -2411
rect 9219 -2501 9225 -2449
rect 11713 -2501 11961 -2449
rect 14449 -2501 15200 -2449
rect 9219 -2539 15200 -2501
rect 15000 -3700 15200 -2539
rect 14994 -3900 15000 -3700
rect 15200 -3900 15206 -3700
rect 14900 -4200 15800 -4000
rect 16000 -4200 16006 -4000
rect 9068 -4238 9132 -4232
rect 9068 -4482 9074 -4238
rect 9126 -4482 9132 -4238
rect 14542 -4238 14606 -4232
rect 9068 -4556 9132 -4482
rect 11805 -4250 11869 -4244
rect 11805 -4494 11811 -4250
rect 11863 -4494 11869 -4250
rect 11805 -4556 11869 -4494
rect 14542 -4482 14548 -4238
rect 14600 -4482 14606 -4238
rect 14542 -4556 14606 -4482
rect 14900 -4556 15100 -4200
rect 15180 -4300 15420 -4280
rect 15180 -4500 15200 -4300
rect 15400 -4500 15800 -4300
rect 16000 -4500 16006 -4300
rect 15180 -4520 15420 -4500
rect 9068 -4620 15100 -4556
rect 12100 -5800 12300 -5794
rect 13600 -5800 13770 -4620
rect 14877 -4899 15117 -4878
rect 14877 -5099 14900 -4899
rect 15100 -5099 15117 -4899
rect 14877 -5122 15117 -5099
rect 9522 -6348 9588 -6341
rect 9522 -6400 9529 -6348
rect 9581 -6400 9588 -6348
rect 9522 -6750 9588 -6400
rect 11650 -6347 11716 -6341
rect 11650 -6399 11657 -6347
rect 11709 -6399 11716 -6347
rect 11650 -6750 11716 -6399
rect 9522 -6810 11716 -6750
rect 10756 -7044 10820 -7038
rect 10756 -7096 10762 -7044
rect 10814 -7096 10820 -7044
rect 10480 -7344 10544 -7338
rect 10480 -7396 10486 -7344
rect 10538 -7396 10544 -7344
rect 10204 -7644 10268 -7638
rect 10204 -7696 10210 -7644
rect 10262 -7696 10268 -7644
rect 9929 -7944 9993 -7938
rect 9929 -7996 9935 -7944
rect 9987 -7996 9993 -7944
rect 9652 -8104 9716 -8100
rect 9652 -8156 9658 -8104
rect 9710 -8156 9716 -8104
rect 9652 -8588 9716 -8156
rect 9652 -8640 9658 -8588
rect 9710 -8640 9716 -8588
rect 9652 -8646 9716 -8640
rect 9929 -8589 9993 -7996
rect 9929 -8641 9935 -8589
rect 9987 -8641 9993 -8589
rect 9929 -8647 9993 -8641
rect 10204 -8588 10268 -7696
rect 10204 -8640 10210 -8588
rect 10262 -8640 10268 -8588
rect 10204 -8646 10268 -8640
rect 10480 -8588 10544 -7396
rect 10480 -8640 10486 -8588
rect 10538 -8640 10544 -8588
rect 10480 -8646 10544 -8640
rect 10756 -8588 10820 -7096
rect 10938 -8390 11002 -6810
rect 10938 -8442 10944 -8390
rect 10996 -8442 11002 -8390
rect 10938 -8448 11002 -8442
rect 10756 -8640 10762 -8588
rect 10814 -8640 10820 -8588
rect 10756 -8646 10820 -8640
rect 9835 -8718 9899 -8712
rect 9835 -8770 9841 -8718
rect 9893 -8770 9899 -8718
rect 9835 -8783 9899 -8770
rect 10111 -8718 10175 -8712
rect 10111 -8770 10117 -8718
rect 10169 -8770 10175 -8718
rect 9835 -8920 9900 -8783
rect 9000 -8980 9900 -8920
rect 10111 -8834 10175 -8770
rect 10387 -8718 10451 -8712
rect 10387 -8770 10393 -8718
rect 10445 -8770 10451 -8718
rect 10111 -8940 10180 -8834
rect 10111 -8942 10182 -8940
rect 10118 -8946 10182 -8942
rect 9000 -19369 9060 -8980
rect 10118 -8998 10124 -8946
rect 10176 -8998 10182 -8946
rect 10118 -9004 10182 -8998
rect 10387 -9040 10451 -8770
rect 10663 -8718 10727 -8712
rect 10663 -8770 10669 -8718
rect 10721 -8770 10727 -8718
rect 10663 -8918 10727 -8770
rect 10663 -9039 10730 -8918
rect 9120 -9100 10451 -9040
rect 10670 -9100 10730 -9039
rect 9120 -17470 9180 -9100
rect 10664 -9160 10670 -9100
rect 10730 -9160 10736 -9100
rect 12100 -9500 12300 -6000
rect 12468 -6000 13770 -5800
rect 12468 -6214 12532 -6000
rect 12468 -8194 12474 -6214
rect 12526 -8194 12532 -6214
rect 12468 -8200 12532 -8194
rect 13706 -6214 13770 -6000
rect 13706 -8194 13712 -6214
rect 13764 -8194 13770 -6214
rect 13706 -8200 13770 -8194
rect 14900 -7800 15100 -5122
rect 15180 -5400 15420 -5380
rect 15780 -5400 16020 -5380
rect 15180 -5600 15200 -5400
rect 15400 -5600 15800 -5400
rect 16000 -5600 16020 -5400
rect 15180 -5620 15420 -5600
rect 15780 -5620 16020 -5600
rect 14580 -8600 14820 -8580
rect 14580 -8800 14600 -8600
rect 14800 -8800 14820 -8600
rect 14580 -8820 14820 -8800
rect 12100 -9706 12300 -9700
rect 14280 -9500 14520 -9480
rect 14280 -9700 14300 -9500
rect 14500 -9700 14520 -9500
rect 14280 -9720 14520 -9700
rect 14300 -12700 14500 -9720
rect 14300 -12906 14500 -12900
rect 14600 -12700 14800 -8820
rect 14600 -12906 14800 -12900
rect 14900 -12700 15100 -8000
rect 15180 -8300 15420 -8280
rect 15180 -8500 15200 -8300
rect 15400 -8500 15420 -8300
rect 15180 -8520 15420 -8500
rect 15200 -9800 15400 -8520
rect 19000 -8700 19200 -8694
rect 15200 -10006 15400 -10000
rect 18700 -9800 18900 -9794
rect 17880 -10400 18120 -10380
rect 17880 -10600 17900 -10400
rect 18100 -10600 18120 -10400
rect 17880 -10620 18120 -10600
rect 17900 -11300 18100 -10620
rect 17900 -11506 18100 -11500
rect 18700 -11200 18900 -10000
rect 19000 -9800 19200 -8900
rect 21100 -9101 21300 -9095
rect 19578 -9500 19816 -9482
rect 19578 -9700 19600 -9500
rect 19800 -9700 19816 -9500
rect 19578 -9721 19816 -9700
rect 19000 -10006 19200 -10000
rect 19600 -11200 19800 -9721
rect 20500 -10100 20700 -10094
rect 20500 -11200 20700 -10300
rect 21100 -11100 21300 -9301
rect 18700 -11300 19100 -11200
rect 18700 -11500 18800 -11300
rect 19000 -11500 19100 -11300
rect 18700 -11600 19100 -11500
rect 19500 -11300 19900 -11200
rect 19500 -11500 19600 -11300
rect 19800 -11500 19900 -11300
rect 19500 -11600 19900 -11500
rect 20400 -11300 20800 -11200
rect 20400 -11500 20500 -11300
rect 20700 -11500 20800 -11300
rect 21100 -11306 21300 -11300
rect 20400 -11600 20800 -11500
rect 14900 -12906 15100 -12900
rect 9280 -17400 9520 -17380
rect 9280 -17470 9300 -17400
rect 9120 -17530 9300 -17470
rect 9280 -17600 9300 -17530
rect 9500 -17600 9520 -17400
rect 9280 -17620 9520 -17600
rect 9280 -19300 9520 -19280
rect 9280 -19369 9300 -19300
rect 9000 -19429 9300 -19369
rect 9280 -19500 9300 -19429
rect 9500 -19500 9520 -19300
rect 9280 -19520 9520 -19500
use sky130_fd_pr__res_xhigh_po_0p69_E9MCU4  R1
timestamp 1716338467
transform 0 1 11699 -1 0 -10331
box -469 -2399 469 2399
use sky130_fd_pr__res_xhigh_po_0p69_39QBTQ  R2
timestamp 1716338467
transform 0 1 16942 -1 0 -11365
box -235 -1442 235 1442
use sky130_fd_pr__res_xhigh_po_0p69_NB3ZKH  R3
timestamp 1716338467
transform 0 1 11745 -1 0 -11414
box -586 -2445 586 2445
use sky130_fd_pr__res_xhigh_po_0p69_GAZAU4  R4
timestamp 1716338467
transform 0 -1 11772 1 0 -13744
box -1756 -2472 1756 2472
use sky130_fd_sc_hd__buf_1  sky130_fd_sc_hd__buf_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 10742 0 1 -8852
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  sky130_fd_sc_hd__buf_1_1
timestamp 1707688321
transform 1 0 9638 0 1 -8852
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  sky130_fd_sc_hd__buf_1_2
timestamp 1707688321
transform 1 0 9914 0 1 -8852
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  sky130_fd_sc_hd__buf_1_3
timestamp 1707688321
transform 1 0 10190 0 1 -8852
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  sky130_fd_sc_hd__buf_1_4
timestamp 1707688321
transform 1 0 10466 0 1 -8852
box -38 -48 314 592
use sbvfcm  x1
timestamp 1716338467
transform 1 0 10300 0 1 -5200
box 5700 -3700 11200 5000
use output_amp  x2
timestamp 1716338467
transform 1 0 10400 0 -1 -14608
box 5100 -2900 11120 4900
use trim_res  x3
timestamp 1716338467
transform 1 0 8600 0 1 -15600
box 700 -3900 5534 -100
use sky130_fd_pr__nfet_01v8_2333C8  XM1
timestamp 1716338467
transform 1 0 11296 0 1 -5340
box -2196 -460 2196 460
use sky130_fd_pr__nfet_01v8_QXBCRM  XM2
timestamp 1716338467
transform 0 -1 14310 1 0 -6704
box -1196 -310 1196 310
use sky130_fd_pr__pfet_01v8_6H4ZLK  XM3
timestamp 1716338467
transform 0 1 13119 -1 0 -7204
box -1196 -719 1196 719
use sky130_fd_pr__pfet_01v8_B3G3L7  XM9
timestamp 1716338467
transform 0 -1 11837 1 0 -2475
box -2225 -2837 2225 2837
use sky130_fd_pr__pfet_01v8_XPMKX6  XM20
timestamp 1716338467
transform 0 1 10619 -1 0 -6374
box -226 -1219 226 1219
<< labels >>
flabel metal1 21300 -10300 21500 -10100 0 FreeSans 256 0 0 0 vbg
port 0 nsew
flabel metal1 21300 -10600 21500 -10400 0 FreeSans 256 0 0 0 vbgtg
port 7 nsew
flabel metal1 21300 -10900 21500 -10700 0 FreeSans 256 0 0 0 vbgsc
port 6 nsew
flabel metal1 21300 -10000 21500 -9800 0 FreeSans 256 0 0 0 vptat
port 13 nsew
flabel metal1 21300 -9700 21500 -9500 0 FreeSans 256 0 0 0 avss
port 1 nsew
flabel metal1 9000 -8600 9200 -8400 0 FreeSans 256 0 0 0 dvdd
port 3 nsew
flabel metal1 9000 -8300 9200 -8100 0 FreeSans 256 0 0 0 trim3
port 8 nsew
flabel metal1 9000 -8000 9200 -7800 0 FreeSans 256 0 0 0 trim2
port 9 nsew
flabel metal1 9000 -7700 9200 -7500 0 FreeSans 256 0 0 0 trim1
port 10 nsew
flabel metal1 9000 -7400 9200 -7200 0 FreeSans 256 0 0 0 trim0
port 11 nsew
flabel metal1 9000 -7100 9200 -6900 0 FreeSans 256 0 0 0 ena
port 5 nsew
flabel metal1 9000 -8900 9200 -8700 0 FreeSans 256 0 0 0 dvss
port 4 nsew
rlabel via1 14900 -8000 15100 -7800 1 vref
flabel metal1 9000 -6600 9200 -6400 0 FreeSans 256 0 0 0 avdd18
port 2 nsew
rlabel metal2 9640 -8980 9700 -8920 1 trim3buf
rlabel metal1 9640 -9040 9700 -8980 1 trim2buf
rlabel metal2 9640 -9100 9700 -9040 1 trim1buf
rlabel metal1 9640 -9160 9700 -9100 1 trim0buf
rlabel metal2 10940 -8240 11000 -8180 1 enabuf
rlabel metal1 9619 -6500 11619 -6456 1 avdd_ena
rlabel via1 15800 -4200 16000 -4000 1 pbias
<< end >>
