magic
tech sky130A
magscale 1 2
timestamp 1719454661
<< ndiff >>
rect 7138 -2690 7196 -1690
rect 8054 -2690 8112 -1690
<< locali >>
rect 6500 4494 6936 4500
rect 6500 4306 6606 4494
rect 6794 4306 6936 4494
rect 6500 4300 6936 4306
<< viali >>
rect 6606 4306 6794 4494
rect 8636 538 8670 4613
rect 10980 532 11014 4607
<< metal1 >>
rect 8380 4880 8620 4900
rect 5319 4748 8119 4876
rect 5168 2644 5232 4692
rect 6406 2650 6470 4692
rect 6600 4520 6800 4748
rect 6580 4494 6820 4520
rect 6580 4306 6606 4494
rect 6794 4306 6820 4494
rect 6580 4280 6820 4306
rect 6400 2644 6476 2650
rect 5168 2580 6406 2644
rect 6470 2580 6476 2644
rect 5700 2520 5900 2580
rect 6400 2574 6476 2580
rect 5680 2500 5920 2520
rect 5680 2300 5700 2500
rect 5900 2300 5920 2500
rect 5680 2280 5920 2300
rect 6600 2200 6800 4280
rect 6968 2650 7032 4692
rect 8206 2650 8270 4692
rect 8380 4680 8400 4880
rect 8600 4834 8620 4880
rect 8600 4706 10850 4834
rect 8600 4680 8620 4706
rect 8380 4660 8620 4680
rect 8616 4613 8744 4619
rect 6962 2644 7038 2650
rect 8200 2644 8276 2650
rect 6962 2580 6968 2644
rect 7032 2580 7038 2644
rect 7119 2580 8119 2644
rect 8200 2580 8206 2644
rect 8270 2580 8276 2644
rect 6962 2574 7038 2580
rect 7500 2520 7700 2580
rect 8200 2574 8276 2580
rect 7480 2500 7720 2520
rect 7480 2300 7500 2500
rect 7700 2300 7720 2500
rect 7480 2280 7720 2300
rect 8616 2200 8636 4613
rect 5100 2000 8636 2200
rect 5100 1700 7000 1900
rect 5100 1400 6700 1600
rect 6500 1194 6700 1400
rect 5328 1130 6700 1194
rect 5267 1052 5331 1058
rect 5267 -936 5273 1052
rect 5325 -936 5331 1052
rect 5267 -942 5331 -936
rect 5725 1052 5789 1058
rect 5725 -493 5731 1052
rect 5783 -493 5789 1052
rect 5725 -942 5789 -493
rect 6183 1052 6247 1058
rect 6183 -936 6189 1052
rect 6241 -936 6247 1052
rect 6183 -942 6247 -936
rect 6500 -1020 6700 1130
rect 5332 -1084 6700 -1020
rect 6500 -1548 6700 -1084
rect 5300 -1612 6700 -1548
rect 5235 -1696 5299 -1690
rect 5235 -2684 5241 -1696
rect 5293 -2684 5299 -1696
rect 5235 -2690 5299 -2684
rect 5693 -1696 5757 -1690
rect 5693 -2294 5699 -1696
rect 5751 -2294 5757 -1696
rect 5693 -2690 5757 -2294
rect 6151 -1696 6215 -1690
rect 6151 -2684 6157 -1696
rect 6209 -2684 6215 -1696
rect 6151 -2690 6215 -2684
rect 6500 -2768 6700 -1612
rect 5300 -2832 6700 -2768
rect 6800 1200 7000 1700
rect 6800 1100 8086 1200
rect 6800 -1020 7000 1100
rect 7167 1052 7231 1058
rect 7167 -936 7173 1052
rect 7225 -936 7231 1052
rect 7167 -942 7231 -936
rect 7625 1052 7689 1058
rect 7625 -494 7631 1052
rect 7683 -494 7689 1052
rect 7625 -942 7689 -494
rect 8083 1052 8147 1058
rect 8083 -936 8089 1052
rect 8141 -936 8147 1052
rect 8500 538 8636 2000
rect 8670 619 8744 4613
rect 9729 1494 9921 4619
rect 9729 625 9735 1494
rect 9915 625 9921 1494
rect 9729 619 9921 625
rect 10906 4607 11034 4619
rect 8670 538 8700 619
rect 8500 300 8700 538
rect 10906 532 10980 4607
rect 11014 532 11034 4607
rect 8800 526 10850 532
rect 8800 410 8806 526
rect 8922 410 10850 526
rect 8800 404 10850 410
rect 10906 300 11034 532
rect 8500 100 11034 300
rect 10100 0 10300 6
rect 8776 -470 8968 -458
rect 8776 -522 8782 -470
rect 8962 -522 8968 -470
rect 8083 -942 8147 -936
rect 8380 -1000 8620 -980
rect 8656 -1000 8720 -600
rect 7690 -1020 8086 -1014
rect 6800 -1084 8086 -1020
rect 6800 -1548 7000 -1084
rect 8380 -1200 8400 -1000
rect 8600 -1200 8720 -1000
rect 8380 -1220 8620 -1200
rect 6800 -1612 8050 -1548
rect 8656 -1600 8720 -1200
rect 9024 -990 9200 -600
rect 9500 -854 9692 -848
rect 9500 -906 9506 -854
rect 9686 -906 9692 -854
rect 9500 -912 9692 -906
rect 9024 -1600 9444 -990
rect 6800 -2768 7000 -1612
rect 7135 -1696 7199 -1690
rect 7135 -2684 7141 -1696
rect 7193 -2684 7199 -1696
rect 7135 -2690 7199 -2684
rect 7593 -1696 7657 -1690
rect 7593 -2294 7599 -1696
rect 7651 -2294 7657 -1696
rect 7593 -2690 7657 -2294
rect 8051 -1696 8115 -1690
rect 8051 -2684 8057 -1696
rect 8109 -2684 8115 -1696
rect 8776 -1740 8968 -1678
rect 8740 -1760 8980 -1740
rect 8740 -1960 8760 -1760
rect 8960 -1960 8980 -1760
rect 8740 -1980 8980 -1960
rect 8051 -2690 8115 -2684
rect 8400 -2046 8968 -1980
rect 8400 -2124 8713 -2046
rect 9200 -2124 9444 -1600
rect 8400 -2624 8720 -2124
rect 9024 -2590 9444 -2124
rect 9748 -1700 9876 -990
rect 10100 -1700 10300 -200
rect 9748 -1900 10300 -1700
rect 9748 -2590 9876 -1900
rect 9024 -2624 9400 -2590
rect 8400 -2702 8714 -2624
rect 8400 -2766 8968 -2702
rect 8400 -2767 8714 -2766
rect 6800 -2832 8050 -2768
rect 8400 -2900 8600 -2767
rect 9200 -2900 9400 -2624
rect 9500 -2674 9692 -2668
rect 9500 -2726 9506 -2674
rect 9686 -2726 9692 -2674
rect 9500 -2732 9692 -2726
rect 10100 -2900 10300 -1900
<< via1 >>
rect 6406 2580 6470 2644
rect 5700 2300 5900 2500
rect 8400 4680 8600 4880
rect 6968 2580 7032 2644
rect 8206 2580 8270 2644
rect 7500 2300 7700 2500
rect 5273 -936 5325 1052
rect 5731 -493 5783 1052
rect 6189 -936 6241 1052
rect 5241 -2684 5293 -1696
rect 5699 -2294 5751 -1696
rect 6157 -2684 6209 -1696
rect 7173 -936 7225 1052
rect 7631 -494 7683 1052
rect 8089 -936 8141 1052
rect 9735 625 9915 1494
rect 8806 410 8922 526
rect 10100 -200 10300 0
rect 8782 -522 8962 -470
rect 8400 -1200 8600 -1000
rect 9506 -906 9686 -854
rect 7141 -2684 7193 -1696
rect 7599 -2294 7651 -1696
rect 8057 -2684 8109 -1696
rect 8760 -1960 8960 -1760
rect 9506 -2726 9686 -2674
<< metal2 >>
rect 8380 4880 8620 4900
rect 8380 4680 8400 4880
rect 8600 4680 8620 4880
rect 8380 4660 8620 4680
rect 6400 2644 6476 2650
rect 6962 2644 7038 2650
rect 8200 2644 8276 2650
rect 6400 2580 6406 2644
rect 6470 2580 6968 2644
rect 7032 2580 8206 2644
rect 8270 2580 8276 2644
rect 6400 2574 6476 2580
rect 6962 2574 7038 2580
rect 8200 2574 8276 2580
rect 5680 2500 5920 2520
rect 5680 2300 5700 2500
rect 5900 2300 5920 2500
rect 5680 2280 5920 2300
rect 7480 2500 7720 2520
rect 8400 2500 8600 4660
rect 7480 2300 7500 2500
rect 7700 2300 8600 2500
rect 7480 2280 7720 2300
rect 5700 1300 5900 2280
rect 7500 1300 7700 2280
rect 5267 1052 5331 1058
rect 5267 -936 5273 1052
rect 5325 -936 5331 1052
rect 5725 1052 5789 1300
rect 5725 -493 5731 1052
rect 5783 -493 5789 1052
rect 5725 -500 5789 -493
rect 6183 1052 6247 1058
rect 5267 -1200 5331 -936
rect 6183 -936 6189 1052
rect 6241 -936 6247 1052
rect 6183 -1200 6247 -936
rect 5267 -1400 6247 -1200
rect 7167 1052 7231 1058
rect 7167 -936 7173 1052
rect 7225 -936 7231 1052
rect 7625 1052 7689 1300
rect 7625 -494 7631 1052
rect 7683 -494 7689 1052
rect 7625 -500 7689 -494
rect 8083 1052 8147 1058
rect 7167 -1200 7231 -936
rect 8083 -936 8089 1052
rect 8141 -936 8147 1052
rect 8300 532 8500 2300
rect 9729 1494 9921 1500
rect 9729 625 9735 1494
rect 9915 625 9921 1494
rect 8300 526 8928 532
rect 8300 410 8806 526
rect 8922 410 8928 526
rect 8300 404 8928 410
rect 8300 0 8500 404
rect 8980 0 9220 20
rect 8300 -200 9000 0
rect 9200 -200 9220 0
rect 9729 0 9921 625
rect 10900 0 11140 20
rect 9729 -200 10100 0
rect 10300 -200 10920 0
rect 11120 -200 11140 0
rect 8980 -220 9220 -200
rect 10900 -220 11140 -200
rect 8776 -470 9200 -458
rect 8776 -522 8782 -470
rect 8962 -522 9200 -470
rect 8776 -528 9200 -522
rect 8083 -1200 8147 -936
rect 9100 -848 9200 -528
rect 9100 -854 9692 -848
rect 9100 -906 9506 -854
rect 9686 -906 9692 -854
rect 9100 -912 9692 -906
rect 7167 -1400 8147 -1200
rect 8380 -1000 8620 -980
rect 8380 -1200 8400 -1000
rect 8600 -1200 8620 -1000
rect 8380 -1220 8620 -1200
rect 5235 -1696 5299 -1690
rect 5235 -2684 5241 -1696
rect 5293 -2400 5299 -1696
rect 5661 -1696 5789 -1400
rect 5661 -2294 5699 -1696
rect 5751 -2294 5789 -1696
rect 5661 -2300 5789 -2294
rect 6151 -1696 6215 -1690
rect 6151 -2400 6157 -1696
rect 5293 -2600 6157 -2400
rect 5293 -2684 5299 -2600
rect 5235 -2690 5299 -2684
rect 6151 -2684 6157 -2600
rect 6209 -2400 6215 -1696
rect 7135 -1696 7199 -1690
rect 7135 -2400 7141 -1696
rect 6209 -2600 7141 -2400
rect 6209 -2684 6215 -2600
rect 6151 -2690 6215 -2684
rect 7135 -2684 7141 -2600
rect 7193 -2400 7199 -1696
rect 7561 -1696 7689 -1400
rect 8400 -1500 8600 -1220
rect 8100 -1690 8600 -1500
rect 7561 -2294 7599 -1696
rect 7651 -2294 7689 -1696
rect 7561 -2300 7689 -2294
rect 8051 -1696 8600 -1690
rect 8051 -2400 8057 -1696
rect 7193 -2600 8057 -2400
rect 7193 -2684 7199 -2600
rect 7135 -2690 7199 -2684
rect 8051 -2684 8057 -2600
rect 8109 -1700 8600 -1696
rect 8109 -2600 8300 -1700
rect 8740 -1760 8980 -1740
rect 8740 -1960 8760 -1760
rect 8960 -1800 8980 -1760
rect 9100 -1800 9200 -912
rect 8960 -1900 9200 -1800
rect 8960 -1960 8980 -1900
rect 8740 -1980 8980 -1960
rect 8109 -2684 8115 -2600
rect 8051 -2690 8115 -2684
rect 9100 -2668 9200 -1900
rect 9100 -2674 9692 -2668
rect 9100 -2726 9506 -2674
rect 9686 -2726 9692 -2674
rect 9100 -2732 9692 -2726
<< via2 >>
rect 9000 -200 9200 0
rect 10920 -200 11120 0
<< metal3 >>
rect 8980 5 9220 20
rect 8980 -205 8995 5
rect 9205 -205 9220 5
rect 8980 -220 9220 -205
rect 10900 5 11140 20
rect 10900 -205 10915 5
rect 11125 -205 11140 5
rect 10900 -220 11140 -205
<< via3 >>
rect 8995 0 9205 5
rect 8995 -200 9000 0
rect 9000 -200 9200 0
rect 9200 -200 9205 0
rect 8995 -205 9205 -200
rect 10915 0 11125 5
rect 10915 -200 10920 0
rect 10920 -200 11120 0
rect 11120 -200 11125 0
rect 10915 -205 11125 -200
<< metal4 >>
rect 8980 5 9220 20
rect 8980 -205 8995 5
rect 9205 0 9220 5
rect 9628 0 10633 345
rect 10900 5 11140 20
rect 10900 0 10915 5
rect 9205 -200 9400 0
rect 9628 -200 10915 0
rect 9205 -205 9220 -200
rect 8980 -220 9220 -205
rect 9628 -658 10633 -200
rect 10900 -205 10915 -200
rect 11125 -205 11140 5
rect 10900 -220 11140 -205
use sky130_fd_pr__cap_mim_m3_1_VCAG9S  XC2
timestamp 1713045697
transform -1 0 9986 0 -1 -160
box -686 -540 686 540
use sky130_fd_pr__nfet_01v8_QGMQL3  XM1
timestamp 1713045697
transform 1 0 8872 0 1 -2374
box -296 -460 296 460
use sky130_fd_pr__nfet_01v8_MMMA4V  XM2
timestamp 1713045697
transform 1 0 8872 0 1 -1100
box -296 -710 296 710
use sky130_fd_pr__nfet_01v8_HS3BL4  XM3
timestamp 1713045697
transform 1 0 9596 0 1 -1790
box -296 -1010 296 1010
use sky130_fd_pr__nfet_01v8_W2FWA4  XM4
timestamp 1713050122
transform 1 0 5725 0 1 -2190
box -625 -710 625 710
use sky130_fd_pr__nfet_01v8_J222PV  XM5
timestamp 1713050122
transform 1 0 7625 0 1 -2190
box -625 -710 625 710
use sky130_fd_pr__pfet_01v8_6H4ZLK  XM6
timestamp 1716081177
transform 0 -1 5819 1 0 3696
box -1196 -719 1196 719
use sky130_fd_pr__pfet_01v8_6H4ZLK  XM7
timestamp 1716081177
transform 0 1 7619 -1 0 3696
box -1196 -719 1196 719
use sky130_fd_pr__pfet_01v8_ST5LSM  XM8
timestamp 1716081120
transform 1 0 9825 0 1 2619
box -1225 -2219 1225 2219
use sky130_fd_pr__nfet_05v0_nvt_CXW7PW  XM9
timestamp 1713050122
transform -1 0 5757 0 -1 58
box -657 -1258 657 1258
use sky130_fd_pr__nfet_05v0_nvt_CXW7PW  XM10
timestamp 1713050122
transform 1 0 7657 0 1 58
box -657 -1258 657 1258
<< labels >>
flabel metal1 5100 1400 5300 1600 0 FreeSans 256 0 0 0 vn
port 3 nsew
flabel metal1 5100 1700 5300 1900 0 FreeSans 256 0 0 0 vp
port 2 nsew
flabel metal1 9200 -2900 9400 -2700 0 FreeSans 256 0 0 0 vss
port 5 nsew
flabel metal1 5100 2000 5300 2200 0 FreeSans 256 0 0 0 vdd
port 0 nsew
flabel metal1 10100 -2900 10300 -2700 0 FreeSans 256 0 0 0 vo
port 1 nsew
flabel metal1 8400 -2900 8600 -2700 0 FreeSans 256 0 0 0 ibias
port 4 nsew
rlabel metal2 8400 -1700 8600 -1500 1 vcm
rlabel via1 7500 2300 7700 2500 1 vo_pre
<< end >>
