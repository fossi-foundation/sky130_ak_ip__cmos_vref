magic
tech sky130A
magscale 1 2
timestamp 1713051387
<< pwell >>
rect -201 -932 201 932
<< psubdiff >>
rect -165 862 -69 896
rect 69 862 165 896
rect -165 800 -131 862
rect 131 800 165 862
rect -165 -862 -131 -800
rect 131 -862 165 -800
rect -165 -896 -69 -862
rect 69 -896 165 -862
<< psubdiffcont >>
rect -69 862 69 896
rect -165 -800 -131 800
rect 131 -800 165 800
rect -69 -896 69 -862
<< xpolycontact >>
rect -35 334 35 766
rect -35 -766 35 -334
<< xpolyres >>
rect -35 -334 35 334
<< locali >>
rect -165 862 -69 896
rect 69 862 165 896
rect -165 800 -131 862
rect 131 800 165 862
rect -165 -862 -131 -800
rect 131 -862 165 -800
rect -165 -896 -69 -862
rect 69 -896 165 -862
<< viali >>
rect -19 351 19 748
rect -19 -748 19 -351
<< metal1 >>
rect -25 748 25 760
rect -25 351 -19 748
rect 19 351 25 748
rect -25 339 25 351
rect -25 -351 25 -339
rect -25 -748 -19 -351
rect 19 -748 25 -351
rect -25 -760 25 -748
<< properties >>
string FIXED_BBOX -148 -879 148 879
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 3.5 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 21.075k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
