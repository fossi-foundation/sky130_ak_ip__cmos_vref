magic
tech sky130A
magscale 1 2
timestamp 1713367752
<< error_p >>
rect 21300 -1594 21320 -1588
rect 21272 -1622 21292 -1616
rect 21274 -4500 21300 -4288
rect 21302 -4528 21328 -4260
rect 20500 -14708 20506 -14702
rect 20694 -14708 20700 -14702
rect 20494 -14714 20500 -14708
rect 20700 -14714 20706 -14708
rect 20494 -14908 20500 -14902
rect 20700 -14908 20706 -14902
rect 20500 -14914 20506 -14908
rect 20694 -14914 20700 -14908
<< error_s >>
rect 16372 -1594 16400 -1588
rect 16400 -1622 16428 -1616
rect 17300 -2194 17306 -2188
rect 17294 -2200 17300 -2194
rect 17294 -2394 17300 -2388
rect 17500 -2394 17506 -2388
rect 9300 -2400 9306 -2394
rect 9494 -2400 9500 -2394
rect 17300 -2400 17306 -2394
rect 17494 -2400 17500 -2394
rect 9294 -2406 9300 -2400
rect 9500 -2406 9506 -2400
rect 9294 -2600 9300 -2594
rect 9500 -2600 9506 -2594
rect 9300 -2606 9306 -2600
rect 9494 -2606 9500 -2600
rect 15462 -3377 15527 -3372
rect 14700 -3400 14706 -3394
rect 14694 -3406 14700 -3400
rect 15434 -3405 15555 -3400
rect 17300 -3494 17306 -3488
rect 17294 -3500 17300 -3494
rect 14694 -3600 14700 -3594
rect 14900 -3600 14906 -3594
rect 14700 -3606 14706 -3600
rect 14894 -3606 14900 -3600
rect 17294 -3694 17300 -3688
rect 17300 -3700 17306 -3694
rect 9300 -4400 9306 -4394
rect 9494 -4400 9500 -4394
rect 9294 -4406 9300 -4400
rect 9500 -4406 9506 -4400
rect 9294 -4600 9300 -4594
rect 9500 -4600 9506 -4594
rect 9300 -4606 9306 -4600
rect 9494 -4606 9500 -4600
rect 18400 -4694 18420 -4688
rect 19272 -4694 19300 -4688
rect 18372 -4722 18392 -4716
rect 19300 -4722 19328 -4716
rect 19200 -5094 19206 -5088
rect 19394 -5094 19400 -5088
rect 19194 -5100 19200 -5094
rect 19400 -5100 19406 -5094
rect 19194 -5294 19200 -5288
rect 19400 -5294 19406 -5288
rect 19200 -5300 19206 -5294
rect 19394 -5300 19400 -5294
rect 19100 -5594 19106 -5588
rect 19294 -5594 19300 -5588
rect 19094 -5600 19100 -5594
rect 19300 -5600 19306 -5594
rect 19094 -5794 19100 -5788
rect 19100 -5800 19106 -5794
rect 14489 -5908 14515 -5903
rect 19472 -6194 19500 -6188
rect 19500 -6222 19528 -6216
rect 18100 -6694 18106 -6688
rect 18294 -6694 18300 -6688
rect 18094 -6700 18100 -6694
rect 18300 -6700 18306 -6694
rect 18094 -6894 18100 -6888
rect 18300 -6894 18306 -6888
rect 18100 -6900 18106 -6894
rect 18294 -6900 18300 -6894
rect 18100 -7694 18106 -7688
rect 18294 -7694 18300 -7688
rect 18094 -7700 18100 -7694
rect 18300 -7700 18306 -7694
rect 18094 -7894 18100 -7888
rect 18300 -7894 18306 -7888
rect 18100 -7900 18106 -7894
rect 18294 -7900 18300 -7894
rect 19400 -9194 19406 -9188
rect 19594 -9194 19600 -9188
rect 19394 -9200 19400 -9194
rect 19600 -9200 19606 -9194
rect 19394 -9394 19400 -9388
rect 19600 -9394 19606 -9388
rect 19400 -9400 19406 -9394
rect 19594 -9400 19600 -9394
rect 19600 -9500 19606 -9494
rect 19794 -9500 19800 -9494
rect 19594 -9506 19600 -9500
rect 19800 -9506 19806 -9500
rect 17900 -10400 17906 -10394
rect 18094 -10400 18100 -10394
rect 17894 -10406 17900 -10400
rect 18100 -10406 18106 -10400
rect 14900 -11700 14906 -11694
rect 15094 -11700 15100 -11694
rect 14894 -11706 14900 -11700
rect 15100 -11706 15106 -11700
rect 19600 -11708 19606 -11702
rect 19794 -11708 19800 -11702
rect 20500 -11708 20506 -11702
rect 20694 -11708 20700 -11702
rect 19594 -11714 19600 -11708
rect 19800 -11714 19806 -11708
rect 20494 -11714 20500 -11708
rect 20700 -11714 20706 -11708
rect 14894 -11900 14900 -11894
rect 15100 -11900 15106 -11894
rect 14900 -11906 14906 -11900
rect 15094 -11906 15100 -11900
rect 19594 -11908 19600 -11902
rect 19800 -11908 19806 -11902
rect 20494 -11908 20500 -11902
rect 20700 -11908 20706 -11902
rect 19600 -11914 19606 -11908
rect 19794 -11914 19800 -11908
rect 20500 -11914 20506 -11908
rect 20694 -11914 20700 -11908
rect 17500 -12008 17506 -12002
rect 17694 -12008 17700 -12002
rect 17494 -12014 17500 -12008
rect 17700 -12014 17706 -12008
rect 17494 -12208 17500 -12202
rect 17700 -12208 17706 -12202
rect 17500 -12214 17506 -12208
rect 17694 -12214 17700 -12208
rect 19000 -13408 19006 -13402
rect 19194 -13408 19200 -13402
rect 18994 -13414 19000 -13408
rect 19200 -13414 19206 -13408
rect 18994 -13608 19000 -13602
rect 19200 -13608 19206 -13602
rect 19000 -13614 19006 -13608
rect 19194 -13614 19200 -13608
rect 10980 -16246 10986 -16240
rect 11174 -16246 11180 -16240
rect 10974 -16252 10980 -16246
rect 11180 -16252 11186 -16246
rect 10974 -16446 10980 -16440
rect 11180 -16446 11186 -16440
rect 10980 -16452 10986 -16446
rect 11174 -16452 11180 -16446
rect 14140 -16560 14146 -16554
rect 14334 -16560 14340 -16554
rect 14134 -16566 14140 -16560
rect 14340 -16566 14346 -16560
rect 13140 -16592 13146 -16586
rect 13146 -16598 13152 -16592
rect 14134 -16760 14140 -16755
rect 14340 -16760 14346 -16755
rect 14140 -16766 14146 -16760
rect 14334 -16766 14340 -16760
<< metal1 >>
rect 9300 -400 9500 -394
rect 9300 -606 9500 -600
rect 11400 -400 11600 -394
rect 11400 -606 11600 -600
rect 12100 -400 12300 -394
rect 14194 -600 14200 -400
rect 14400 -600 14406 -400
rect 12100 -606 12300 -600
rect 9100 -1500 14900 -1300
rect 12000 -2400 12200 -2394
rect 11394 -2600 11400 -2400
rect 11600 -2600 11606 -2400
rect 12000 -2606 12200 -2600
rect 14200 -2400 14400 -2394
rect 14200 -2606 14400 -2600
rect 14700 -3400 14900 -1500
rect 15200 -1900 15400 -200
rect 15500 -400 15700 -200
rect 15591 -1172 15660 -400
rect 15465 -1241 15471 -1172
rect 15540 -1241 15660 -1172
rect 15694 -1500 15700 -1300
rect 15900 -1500 15906 -1300
rect 15700 -1894 15900 -1500
rect 15200 -2100 15600 -1900
rect 15700 -2094 16300 -1894
rect 15200 -2103 15400 -2100
rect 9100 -3600 14700 -3400
rect 15000 -2400 15200 -2394
rect 11500 -4400 11700 -4394
rect 11500 -4606 11700 -4600
rect 12000 -4400 12200 -4394
rect 12000 -4606 12200 -4600
rect 14200 -4400 14400 -4394
rect 14200 -4606 14400 -4600
rect 15000 -5000 15200 -2600
rect 15462 -3319 15527 -3313
rect 15462 -3371 15469 -3319
rect 15521 -3322 15527 -3319
rect 15521 -3368 15659 -3322
rect 15521 -3371 15527 -3368
rect 15462 -3377 15527 -3371
rect 8999 -5790 9290 -5289
rect 9400 -5400 13200 -5200
rect 15000 -5206 15200 -5200
rect 15700 -4400 15900 -2094
rect 13000 -5700 13200 -5400
rect 9000 -8900 9200 -5790
rect 9400 -5900 13200 -5700
rect 13302 -5300 13450 -5286
rect 13302 -5500 15200 -5300
rect 15400 -5500 15406 -5300
rect 13302 -5794 13450 -5500
rect 14206 -5898 14414 -5500
rect 13000 -6000 13200 -5900
rect 14487 -5969 14489 -5903
rect 14131 -6000 14489 -5969
rect 12300 -6200 12500 -6194
rect 13000 -6200 14489 -6000
rect 12300 -6700 12500 -6400
rect 12614 -6500 12700 -6300
rect 12900 -6500 13400 -6300
rect 13600 -6500 13623 -6300
rect 12700 -6504 13623 -6500
rect 12300 -6900 13700 -6700
rect 12500 -8400 12700 -6900
rect 13500 -8400 13700 -6900
rect 14131 -7900 14489 -6200
rect 15700 -6300 15900 -4600
rect 16000 -2394 16800 -2194
rect 16000 -3400 16200 -2394
rect 16000 -4700 16200 -3600
rect 15994 -4900 16000 -4700
rect 16200 -4900 16206 -4700
rect 16100 -5000 16300 -4994
rect 16100 -5206 16300 -5200
rect 14594 -6500 14600 -6300
rect 14800 -6500 15900 -6300
rect 14880 -7900 15120 -7880
rect 14131 -8100 14900 -7900
rect 15100 -8100 15120 -7900
rect 14880 -8120 15120 -8100
rect 14300 -8400 15200 -8200
rect 15400 -8400 15406 -8200
rect 12700 -8600 13600 -8500
rect 14300 -8600 14500 -8400
rect 12700 -8800 14500 -8600
rect 14580 -8600 14820 -8580
rect 15700 -8600 15900 -6500
rect 14580 -8800 14600 -8600
rect 14800 -8800 15900 -8600
rect 14580 -8820 14820 -8800
rect 9000 -9100 14300 -8900
rect 14500 -9100 16000 -8900
rect 9172 -9456 13000 -9338
rect 13205 -9456 14800 -9338
rect 12900 -9572 13000 -9456
rect 9172 -9924 9593 -9572
rect 12900 -9690 13626 -9572
rect 13205 -9924 14500 -9806
rect 9172 -10656 9593 -10304
rect 13297 -10422 14200 -10304
rect 9172 -11124 9593 -10772
rect 13297 -10890 13718 -10538
rect 14000 -10700 14200 -10422
rect 14300 -10400 14500 -9924
rect 14600 -10100 14800 -9456
rect 15800 -9500 16000 -9100
rect 19700 -9500 19900 -9194
rect 15800 -9700 19600 -9500
rect 19800 -9700 19900 -9500
rect 15194 -10000 15200 -9800
rect 15400 -10000 18700 -9800
rect 18900 -10000 18906 -9800
rect 20994 -10000 21000 -9800
rect 21200 -10000 21500 -9800
rect 14600 -10300 20500 -10100
rect 20700 -10300 21500 -10100
rect 14300 -10600 17900 -10400
rect 18100 -10600 21500 -10400
rect 14000 -10900 21500 -10700
rect 13297 -11124 14200 -11006
rect 14000 -11464 14200 -11124
rect 15800 -11400 16000 -10900
rect 9172 -11816 9593 -11464
rect 13351 -11582 15400 -11464
rect 17894 -11500 17900 -11300
rect 18100 -11500 18106 -11300
rect 9172 -12284 9593 -11932
rect 13351 -12050 13772 -11698
rect 14300 -11700 14500 -11694
rect 9172 -12752 9593 -12400
rect 13351 -12518 13772 -12166
rect 9172 -13220 9593 -12868
rect 13351 -12986 13772 -12634
rect 9172 -13688 9593 -13336
rect 13351 -13454 13772 -13102
rect 9172 -14156 9593 -13804
rect 13351 -13922 13772 -13570
rect 9172 -14624 9593 -14272
rect 13351 -14390 13772 -14038
rect 11640 -14624 13772 -14506
rect 11640 -15060 11840 -14624
rect 14300 -14860 14500 -11900
rect 11900 -15060 14500 -14860
rect 14600 -11700 14800 -11694
rect 9000 -15300 9200 -15100
rect 9000 -15600 9200 -15400
rect 14600 -16608 14800 -11900
rect 14900 -16308 15100 -11900
rect 15200 -16008 15400 -11582
rect 18700 -11708 18900 -11702
rect 18700 -11914 18900 -11908
rect 15200 -16208 15700 -16008
rect 14900 -16508 15700 -16308
rect 14600 -16808 15700 -16608
rect 9000 -19200 9200 -19000
rect 9000 -19500 9200 -19300
rect 14600 -19500 14800 -19300
rect 15200 -19500 15400 -19300
<< via1 >>
rect 9300 -600 9500 -400
rect 11400 -600 11600 -400
rect 12100 -600 12300 -400
rect 14200 -600 14400 -400
rect 9300 -2600 9500 -2400
rect 11400 -2600 11600 -2400
rect 12000 -2600 12200 -2400
rect 14200 -2600 14400 -2400
rect 15471 -1241 15540 -1172
rect 15700 -1500 15900 -1300
rect 14700 -3600 14900 -3400
rect 15000 -2600 15200 -2400
rect 9300 -4600 9500 -4400
rect 11500 -4600 11700 -4400
rect 12000 -4600 12200 -4400
rect 14200 -4600 14400 -4400
rect 15469 -3371 15521 -3319
rect 15000 -5200 15200 -5000
rect 15700 -4600 15900 -4400
rect 15200 -5500 15400 -5300
rect 12300 -6400 12500 -6200
rect 12700 -6500 12900 -6300
rect 13400 -6500 13600 -6300
rect 16000 -3600 16200 -3400
rect 16000 -4900 16200 -4700
rect 16100 -5200 16300 -5000
rect 14600 -6500 14800 -6300
rect 14900 -8100 15100 -7900
rect 15200 -8400 15400 -8200
rect 14600 -8800 14800 -8600
rect 14300 -9100 14500 -8900
rect 19400 -9394 19600 -9194
rect 19600 -9700 19800 -9500
rect 15200 -10000 15400 -9800
rect 18700 -10000 18900 -9800
rect 21000 -10000 21200 -9800
rect 20500 -10300 20700 -10100
rect 17900 -10600 18100 -10400
rect 17900 -11500 18100 -11300
rect 14300 -11900 14500 -11700
rect 14600 -11900 14800 -11700
rect 14900 -11900 15100 -11700
rect 18700 -11908 18900 -11708
rect 19600 -11908 19800 -11708
rect 20500 -11908 20700 -11708
<< metal2 >>
rect 14200 -400 14400 -394
rect 9294 -600 9300 -400
rect 9500 -600 11400 -400
rect 11600 -600 12100 -400
rect 12300 -600 14200 -400
rect 14200 -800 14400 -600
rect 14200 -1000 15900 -800
rect 15471 -1172 15540 -1166
rect 15471 -1247 15540 -1241
rect 11400 -2400 11600 -2394
rect 9500 -2600 11400 -2400
rect 11600 -2600 12000 -2400
rect 12200 -2600 14200 -2400
rect 14400 -2600 15000 -2400
rect 15200 -2600 15206 -2400
rect 11400 -2606 11600 -2600
rect 15472 -3313 15518 -1247
rect 15700 -1300 15900 -1000
rect 15700 -1506 15900 -1500
rect 15462 -3319 15527 -3313
rect 15462 -3371 15469 -3319
rect 15521 -3371 15527 -3319
rect 15462 -3377 15527 -3371
rect 14900 -3600 16000 -3400
rect 16200 -3600 16206 -3400
rect 9500 -4600 11500 -4400
rect 11700 -4600 12000 -4400
rect 12200 -4600 14200 -4400
rect 14400 -4600 15700 -4400
rect 15900 -4600 15906 -4400
rect 16000 -4700 16200 -4694
rect 12300 -4900 16000 -4700
rect 12300 -6200 12500 -4900
rect 16000 -4906 16200 -4900
rect 14900 -5200 15000 -5000
rect 15200 -5200 16100 -5000
rect 16300 -5200 16306 -5000
rect 12294 -6400 12300 -6200
rect 12500 -6400 12506 -6200
rect 14600 -6300 14800 -6294
rect 12614 -6500 12700 -6300
rect 12900 -6500 13400 -6300
rect 13600 -6500 14600 -6300
rect 12700 -6504 13623 -6500
rect 13400 -6506 13600 -6504
rect 14600 -6506 14800 -6500
rect 14900 -7880 15100 -5200
rect 15200 -5300 15400 -5294
rect 15400 -5500 16700 -5300
rect 15200 -5506 15400 -5500
rect 14880 -7900 15120 -7880
rect 14880 -8100 14900 -7900
rect 15100 -8100 15120 -7900
rect 14880 -8120 15120 -8100
rect 14580 -8600 14820 -8580
rect 14580 -8800 14600 -8600
rect 14800 -8800 14820 -8600
rect 14580 -8820 14820 -8800
rect 14300 -8900 14500 -8893
rect 14300 -11700 14500 -9100
rect 14600 -11700 14800 -8820
rect 14900 -11700 15100 -8120
rect 15200 -8200 15400 -8194
rect 15200 -9800 15400 -8400
rect 19600 -9394 21200 -9194
rect 15200 -10006 15400 -10000
rect 18700 -9800 18900 -9794
rect 17900 -11300 18100 -10600
rect 17900 -11506 18100 -11500
rect 14294 -11900 14300 -11700
rect 14500 -11900 14506 -11700
rect 14594 -11900 14600 -11700
rect 14800 -11900 14806 -11700
rect 18700 -11708 18900 -10000
rect 19600 -11708 19800 -9700
rect 21000 -9800 21200 -9394
rect 21000 -10006 21200 -10000
rect 18694 -11908 18700 -11708
rect 18900 -11908 18906 -11708
rect 20500 -10100 20700 -10094
rect 20500 -11708 20700 -10300
use sky130_fd_pr__res_xhigh_po_0p69_E9MCU4  R1
timestamp 1713140876
transform 0 1 11399 -1 0 -9631
box -469 -2399 469 2399
use sky130_fd_pr__res_xhigh_po_0p69_39QBTQ  R2
timestamp 1713056482
transform 0 1 16942 -1 0 -11365
box -235 -1442 235 1442
use sky130_fd_pr__res_xhigh_po_0p69_NB3ZKH  R3
timestamp 1713140876
transform 0 1 11445 -1 0 -10714
box -586 -2445 586 2445
use sky130_fd_pr__res_xhigh_po_0p69_GAZAU4  R4
timestamp 1713140876
transform 0 -1 11472 1 0 -13044
box -1756 -2472 1756 2472
use sbvfcm  x1
timestamp 1713214705
transform 1 0 10400 0 1 -5694
box 5700 -3706 11200 5500
use output_amp  x2
timestamp 1713362954
transform 1 0 10400 0 -1 -14608
box 5100 -2903 11050 4892
use trim_res  x3
timestamp 1713116496
transform 1 0 8480 0 1 -15320
box 720 -4180 5972 460
use sky130_fd_pr__nfet_01v8_2333C8  XM1
timestamp 1713045697
transform 1 0 11296 0 1 -5540
box -2196 -460 2196 460
use sky130_fd_pr__nfet_01v8_QXBCRM  XM2
timestamp 1713051622
transform 0 -1 14310 1 0 -6904
box -1196 -310 1196 310
use sky130_fd_pr__pfet_01v8_6H4ZLK  XM3
timestamp 1713045697
transform 0 1 13119 -1 0 -7504
box -1196 -719 1196 719
use sky130_fd_pr__pfet_01v8_B3G3L7  XM9
timestamp 1713056482
transform 0 -1 11837 1 0 -2475
box -2225 -2837 2225 2837
use sky130_fd_pr__pfet_01v8_XPMKX6  XM20
timestamp 1713045697
transform 1 0 15626 0 1 -2281
box -226 -1219 226 1219
<< labels >>
flabel metal1 21300 -10300 21500 -10100 0 FreeSans 256 0 0 0 vbg
port 0 nsew
flabel metal1 21300 -10600 21500 -10400 0 FreeSans 256 0 0 0 vbgtg
port 7 nsew
flabel metal1 21300 -10900 21500 -10700 0 FreeSans 256 0 0 0 vbgsc
port 6 nsew
flabel metal1 9000 -19500 9200 -19300 0 FreeSans 256 0 0 0 trim3
port 8 nsew
flabel metal1 9000 -19200 9200 -19000 0 FreeSans 256 0 0 0 trim2
port 9 nsew
flabel metal1 9000 -15600 9200 -15400 0 FreeSans 256 0 0 0 trim0
port 11 nsew
flabel metal1 9000 -15300 9200 -15100 0 FreeSans 256 0 0 0 trim1
port 10 nsew
flabel metal1 9000 -9100 9200 -8900 0 FreeSans 256 0 0 0 avss
port 1 nsew
flabel metal1 21300 -10000 21500 -9800 0 FreeSans 256 0 0 0 vptat
port 13 nsew
flabel metal1 14600 -19500 14800 -19300 0 FreeSans 256 0 0 0 dvdd
port 3 nsew
flabel metal1 15200 -400 15400 -200 0 FreeSans 256 0 0 0 avdd18
port 2 nsew
flabel metal1 15500 -400 15700 -200 0 FreeSans 256 0 0 0 ena
port 5 nsew
flabel metal1 15200 -19500 15400 -19300 0 FreeSans 256 0 0 0 dvss
port 4 nsew
<< end >>
