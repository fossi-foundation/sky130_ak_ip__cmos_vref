magic
tech sky130A
magscale 1 2
timestamp 1713212409
<< pwell >>
rect -3831 -835 3831 835
<< nmos >>
rect -3635 -625 -3235 625
rect -3177 -625 -2777 625
rect -2719 -625 -2319 625
rect -2261 -625 -1861 625
rect -1803 -625 -1403 625
rect -1345 -625 -945 625
rect -887 -625 -487 625
rect -429 -625 -29 625
rect 29 -625 429 625
rect 487 -625 887 625
rect 945 -625 1345 625
rect 1403 -625 1803 625
rect 1861 -625 2261 625
rect 2319 -625 2719 625
rect 2777 -625 3177 625
rect 3235 -625 3635 625
<< ndiff >>
rect -3693 613 -3635 625
rect -3693 -613 -3681 613
rect -3647 -613 -3635 613
rect -3693 -625 -3635 -613
rect -3235 613 -3177 625
rect -3235 -613 -3223 613
rect -3189 -613 -3177 613
rect -3235 -625 -3177 -613
rect -2777 613 -2719 625
rect -2777 -613 -2765 613
rect -2731 -613 -2719 613
rect -2777 -625 -2719 -613
rect -2319 613 -2261 625
rect -2319 -613 -2307 613
rect -2273 -613 -2261 613
rect -2319 -625 -2261 -613
rect -1861 613 -1803 625
rect -1861 -613 -1849 613
rect -1815 -613 -1803 613
rect -1861 -625 -1803 -613
rect -1403 613 -1345 625
rect -1403 -613 -1391 613
rect -1357 -613 -1345 613
rect -1403 -625 -1345 -613
rect -945 613 -887 625
rect -945 -613 -933 613
rect -899 -613 -887 613
rect -945 -625 -887 -613
rect -487 613 -429 625
rect -487 -613 -475 613
rect -441 -613 -429 613
rect -487 -625 -429 -613
rect -29 613 29 625
rect -29 -613 -17 613
rect 17 -613 29 613
rect -29 -625 29 -613
rect 429 613 487 625
rect 429 -613 441 613
rect 475 -613 487 613
rect 429 -625 487 -613
rect 887 613 945 625
rect 887 -613 899 613
rect 933 -613 945 613
rect 887 -625 945 -613
rect 1345 613 1403 625
rect 1345 -613 1357 613
rect 1391 -613 1403 613
rect 1345 -625 1403 -613
rect 1803 613 1861 625
rect 1803 -613 1815 613
rect 1849 -613 1861 613
rect 1803 -625 1861 -613
rect 2261 613 2319 625
rect 2261 -613 2273 613
rect 2307 -613 2319 613
rect 2261 -625 2319 -613
rect 2719 613 2777 625
rect 2719 -613 2731 613
rect 2765 -613 2777 613
rect 2719 -625 2777 -613
rect 3177 613 3235 625
rect 3177 -613 3189 613
rect 3223 -613 3235 613
rect 3177 -625 3235 -613
rect 3635 613 3693 625
rect 3635 -613 3647 613
rect 3681 -613 3693 613
rect 3635 -625 3693 -613
<< ndiffc >>
rect -3681 -613 -3647 613
rect -3223 -613 -3189 613
rect -2765 -613 -2731 613
rect -2307 -613 -2273 613
rect -1849 -613 -1815 613
rect -1391 -613 -1357 613
rect -933 -613 -899 613
rect -475 -613 -441 613
rect -17 -613 17 613
rect 441 -613 475 613
rect 899 -613 933 613
rect 1357 -613 1391 613
rect 1815 -613 1849 613
rect 2273 -613 2307 613
rect 2731 -613 2765 613
rect 3189 -613 3223 613
rect 3647 -613 3681 613
<< psubdiff >>
rect -3795 765 -3699 799
rect 3699 765 3795 799
rect -3795 703 -3761 765
rect 3761 703 3795 765
rect -3795 -765 -3761 -703
rect 3761 -765 3795 -703
rect -3795 -799 -3699 -765
rect 3699 -799 3795 -765
<< psubdiffcont >>
rect -3699 765 3699 799
rect -3795 -703 -3761 703
rect 3761 -703 3795 703
rect -3699 -799 3699 -765
<< poly >>
rect -3635 697 -3235 713
rect -3635 663 -3619 697
rect -3251 663 -3235 697
rect -3635 625 -3235 663
rect -3177 697 -2777 713
rect -3177 663 -3161 697
rect -2793 663 -2777 697
rect -3177 625 -2777 663
rect -2719 697 -2319 713
rect -2719 663 -2703 697
rect -2335 663 -2319 697
rect -2719 625 -2319 663
rect -2261 697 -1861 713
rect -2261 663 -2245 697
rect -1877 663 -1861 697
rect -2261 625 -1861 663
rect -1803 697 -1403 713
rect -1803 663 -1787 697
rect -1419 663 -1403 697
rect -1803 625 -1403 663
rect -1345 697 -945 713
rect -1345 663 -1329 697
rect -961 663 -945 697
rect -1345 625 -945 663
rect -887 697 -487 713
rect -887 663 -871 697
rect -503 663 -487 697
rect -887 625 -487 663
rect -429 697 -29 713
rect -429 663 -413 697
rect -45 663 -29 697
rect -429 625 -29 663
rect 29 697 429 713
rect 29 663 45 697
rect 413 663 429 697
rect 29 625 429 663
rect 487 697 887 713
rect 487 663 503 697
rect 871 663 887 697
rect 487 625 887 663
rect 945 697 1345 713
rect 945 663 961 697
rect 1329 663 1345 697
rect 945 625 1345 663
rect 1403 697 1803 713
rect 1403 663 1419 697
rect 1787 663 1803 697
rect 1403 625 1803 663
rect 1861 697 2261 713
rect 1861 663 1877 697
rect 2245 663 2261 697
rect 1861 625 2261 663
rect 2319 697 2719 713
rect 2319 663 2335 697
rect 2703 663 2719 697
rect 2319 625 2719 663
rect 2777 697 3177 713
rect 2777 663 2793 697
rect 3161 663 3177 697
rect 2777 625 3177 663
rect 3235 697 3635 713
rect 3235 663 3251 697
rect 3619 663 3635 697
rect 3235 625 3635 663
rect -3635 -663 -3235 -625
rect -3635 -697 -3619 -663
rect -3251 -697 -3235 -663
rect -3635 -713 -3235 -697
rect -3177 -663 -2777 -625
rect -3177 -697 -3161 -663
rect -2793 -697 -2777 -663
rect -3177 -713 -2777 -697
rect -2719 -663 -2319 -625
rect -2719 -697 -2703 -663
rect -2335 -697 -2319 -663
rect -2719 -713 -2319 -697
rect -2261 -663 -1861 -625
rect -2261 -697 -2245 -663
rect -1877 -697 -1861 -663
rect -2261 -713 -1861 -697
rect -1803 -663 -1403 -625
rect -1803 -697 -1787 -663
rect -1419 -697 -1403 -663
rect -1803 -713 -1403 -697
rect -1345 -663 -945 -625
rect -1345 -697 -1329 -663
rect -961 -697 -945 -663
rect -1345 -713 -945 -697
rect -887 -663 -487 -625
rect -887 -697 -871 -663
rect -503 -697 -487 -663
rect -887 -713 -487 -697
rect -429 -663 -29 -625
rect -429 -697 -413 -663
rect -45 -697 -29 -663
rect -429 -713 -29 -697
rect 29 -663 429 -625
rect 29 -697 45 -663
rect 413 -697 429 -663
rect 29 -713 429 -697
rect 487 -663 887 -625
rect 487 -697 503 -663
rect 871 -697 887 -663
rect 487 -713 887 -697
rect 945 -663 1345 -625
rect 945 -697 961 -663
rect 1329 -697 1345 -663
rect 945 -713 1345 -697
rect 1403 -663 1803 -625
rect 1403 -697 1419 -663
rect 1787 -697 1803 -663
rect 1403 -713 1803 -697
rect 1861 -663 2261 -625
rect 1861 -697 1877 -663
rect 2245 -697 2261 -663
rect 1861 -713 2261 -697
rect 2319 -663 2719 -625
rect 2319 -697 2335 -663
rect 2703 -697 2719 -663
rect 2319 -713 2719 -697
rect 2777 -663 3177 -625
rect 2777 -697 2793 -663
rect 3161 -697 3177 -663
rect 2777 -713 3177 -697
rect 3235 -663 3635 -625
rect 3235 -697 3251 -663
rect 3619 -697 3635 -663
rect 3235 -713 3635 -697
<< polycont >>
rect -3619 663 -3251 697
rect -3161 663 -2793 697
rect -2703 663 -2335 697
rect -2245 663 -1877 697
rect -1787 663 -1419 697
rect -1329 663 -961 697
rect -871 663 -503 697
rect -413 663 -45 697
rect 45 663 413 697
rect 503 663 871 697
rect 961 663 1329 697
rect 1419 663 1787 697
rect 1877 663 2245 697
rect 2335 663 2703 697
rect 2793 663 3161 697
rect 3251 663 3619 697
rect -3619 -697 -3251 -663
rect -3161 -697 -2793 -663
rect -2703 -697 -2335 -663
rect -2245 -697 -1877 -663
rect -1787 -697 -1419 -663
rect -1329 -697 -961 -663
rect -871 -697 -503 -663
rect -413 -697 -45 -663
rect 45 -697 413 -663
rect 503 -697 871 -663
rect 961 -697 1329 -663
rect 1419 -697 1787 -663
rect 1877 -697 2245 -663
rect 2335 -697 2703 -663
rect 2793 -697 3161 -663
rect 3251 -697 3619 -663
<< locali >>
rect -3795 765 -3699 799
rect 3699 765 3795 799
rect -3795 703 -3761 765
rect 3761 703 3795 765
rect -3635 663 -3619 697
rect -3251 663 -3235 697
rect -3177 663 -3161 697
rect -2793 663 -2777 697
rect -2719 663 -2703 697
rect -2335 663 -2319 697
rect -2261 663 -2245 697
rect -1877 663 -1861 697
rect -1803 663 -1787 697
rect -1419 663 -1403 697
rect -1345 663 -1329 697
rect -961 663 -945 697
rect -887 663 -871 697
rect -503 663 -487 697
rect -429 663 -413 697
rect -45 663 -29 697
rect 29 663 45 697
rect 413 663 429 697
rect 487 663 503 697
rect 871 663 887 697
rect 945 663 961 697
rect 1329 663 1345 697
rect 1403 663 1419 697
rect 1787 663 1803 697
rect 1861 663 1877 697
rect 2245 663 2261 697
rect 2319 663 2335 697
rect 2703 663 2719 697
rect 2777 663 2793 697
rect 3161 663 3177 697
rect 3235 663 3251 697
rect 3619 663 3635 697
rect -3681 613 -3647 629
rect -3681 -629 -3647 -613
rect -3223 613 -3189 629
rect -3223 -629 -3189 -613
rect -2765 613 -2731 629
rect -2765 -629 -2731 -613
rect -2307 613 -2273 629
rect -2307 -629 -2273 -613
rect -1849 613 -1815 629
rect -1849 -629 -1815 -613
rect -1391 613 -1357 629
rect -1391 -629 -1357 -613
rect -933 613 -899 629
rect -933 -629 -899 -613
rect -475 613 -441 629
rect -475 -629 -441 -613
rect -17 613 17 629
rect -17 -629 17 -613
rect 441 613 475 629
rect 441 -629 475 -613
rect 899 613 933 629
rect 899 -629 933 -613
rect 1357 613 1391 629
rect 1357 -629 1391 -613
rect 1815 613 1849 629
rect 1815 -629 1849 -613
rect 2273 613 2307 629
rect 2273 -629 2307 -613
rect 2731 613 2765 629
rect 2731 -629 2765 -613
rect 3189 613 3223 629
rect 3189 -629 3223 -613
rect 3647 613 3681 629
rect 3647 -629 3681 -613
rect -3635 -697 -3619 -663
rect -3251 -697 -3235 -663
rect -3177 -697 -3161 -663
rect -2793 -697 -2777 -663
rect -2719 -697 -2703 -663
rect -2335 -697 -2319 -663
rect -2261 -697 -2245 -663
rect -1877 -697 -1861 -663
rect -1803 -697 -1787 -663
rect -1419 -697 -1403 -663
rect -1345 -697 -1329 -663
rect -961 -697 -945 -663
rect -887 -697 -871 -663
rect -503 -697 -487 -663
rect -429 -697 -413 -663
rect -45 -697 -29 -663
rect 29 -697 45 -663
rect 413 -697 429 -663
rect 487 -697 503 -663
rect 871 -697 887 -663
rect 945 -697 961 -663
rect 1329 -697 1345 -663
rect 1403 -697 1419 -663
rect 1787 -697 1803 -663
rect 1861 -697 1877 -663
rect 2245 -697 2261 -663
rect 2319 -697 2335 -663
rect 2703 -697 2719 -663
rect 2777 -697 2793 -663
rect 3161 -697 3177 -663
rect 3235 -697 3251 -663
rect 3619 -697 3635 -663
rect -3795 -765 -3761 -703
rect 3761 -765 3795 -703
rect -3795 -799 -3699 -765
rect 3699 -799 3795 -765
<< viali >>
rect -3619 663 -3251 697
rect -3161 663 -2793 697
rect -2703 663 -2335 697
rect -2245 663 -1877 697
rect -1787 663 -1419 697
rect -1329 663 -961 697
rect -871 663 -503 697
rect -413 663 -45 697
rect 45 663 413 697
rect 503 663 871 697
rect 961 663 1329 697
rect 1419 663 1787 697
rect 1877 663 2245 697
rect 2335 663 2703 697
rect 2793 663 3161 697
rect 3251 663 3619 697
rect -3681 -613 -3647 613
rect -3223 -613 -3189 613
rect -2765 -613 -2731 613
rect -2307 -613 -2273 613
rect -1849 -613 -1815 613
rect -1391 -613 -1357 613
rect -933 -613 -899 613
rect -475 -613 -441 613
rect -17 -613 17 613
rect 441 -613 475 613
rect 899 -613 933 613
rect 1357 -613 1391 613
rect 1815 -613 1849 613
rect 2273 -613 2307 613
rect 2731 -613 2765 613
rect 3189 -613 3223 613
rect 3647 -613 3681 613
rect -3619 -697 -3251 -663
rect -3161 -697 -2793 -663
rect -2703 -697 -2335 -663
rect -2245 -697 -1877 -663
rect -1787 -697 -1419 -663
rect -1329 -697 -961 -663
rect -871 -697 -503 -663
rect -413 -697 -45 -663
rect 45 -697 413 -663
rect 503 -697 871 -663
rect 961 -697 1329 -663
rect 1419 -697 1787 -663
rect 1877 -697 2245 -663
rect 2335 -697 2703 -663
rect 2793 -697 3161 -663
rect 3251 -697 3619 -663
<< metal1 >>
rect -3631 697 -3239 703
rect -3631 663 -3619 697
rect -3251 663 -3239 697
rect -3631 657 -3239 663
rect -3173 697 -2781 703
rect -3173 663 -3161 697
rect -2793 663 -2781 697
rect -3173 657 -2781 663
rect -2715 697 -2323 703
rect -2715 663 -2703 697
rect -2335 663 -2323 697
rect -2715 657 -2323 663
rect -2257 697 -1865 703
rect -2257 663 -2245 697
rect -1877 663 -1865 697
rect -2257 657 -1865 663
rect -1799 697 -1407 703
rect -1799 663 -1787 697
rect -1419 663 -1407 697
rect -1799 657 -1407 663
rect -1341 697 -949 703
rect -1341 663 -1329 697
rect -961 663 -949 697
rect -1341 657 -949 663
rect -883 697 -491 703
rect -883 663 -871 697
rect -503 663 -491 697
rect -883 657 -491 663
rect -425 697 -33 703
rect -425 663 -413 697
rect -45 663 -33 697
rect -425 657 -33 663
rect 33 697 425 703
rect 33 663 45 697
rect 413 663 425 697
rect 33 657 425 663
rect 491 697 883 703
rect 491 663 503 697
rect 871 663 883 697
rect 491 657 883 663
rect 949 697 1341 703
rect 949 663 961 697
rect 1329 663 1341 697
rect 949 657 1341 663
rect 1407 697 1799 703
rect 1407 663 1419 697
rect 1787 663 1799 697
rect 1407 657 1799 663
rect 1865 697 2257 703
rect 1865 663 1877 697
rect 2245 663 2257 697
rect 1865 657 2257 663
rect 2323 697 2715 703
rect 2323 663 2335 697
rect 2703 663 2715 697
rect 2323 657 2715 663
rect 2781 697 3173 703
rect 2781 663 2793 697
rect 3161 663 3173 697
rect 2781 657 3173 663
rect 3239 697 3631 703
rect 3239 663 3251 697
rect 3619 663 3631 697
rect 3239 657 3631 663
rect -3687 613 -3641 625
rect -3687 -613 -3681 613
rect -3647 -613 -3641 613
rect -3687 -625 -3641 -613
rect -3229 613 -3183 625
rect -3229 -613 -3223 613
rect -3189 -613 -3183 613
rect -3229 -625 -3183 -613
rect -2771 613 -2725 625
rect -2771 -613 -2765 613
rect -2731 -613 -2725 613
rect -2771 -625 -2725 -613
rect -2313 613 -2267 625
rect -2313 -613 -2307 613
rect -2273 -613 -2267 613
rect -2313 -625 -2267 -613
rect -1855 613 -1809 625
rect -1855 -613 -1849 613
rect -1815 -613 -1809 613
rect -1855 -625 -1809 -613
rect -1397 613 -1351 625
rect -1397 -613 -1391 613
rect -1357 -613 -1351 613
rect -1397 -625 -1351 -613
rect -939 613 -893 625
rect -939 -613 -933 613
rect -899 -613 -893 613
rect -939 -625 -893 -613
rect -481 613 -435 625
rect -481 -613 -475 613
rect -441 -613 -435 613
rect -481 -625 -435 -613
rect -23 613 23 625
rect -23 -613 -17 613
rect 17 -613 23 613
rect -23 -625 23 -613
rect 435 613 481 625
rect 435 -613 441 613
rect 475 -613 481 613
rect 435 -625 481 -613
rect 893 613 939 625
rect 893 -613 899 613
rect 933 -613 939 613
rect 893 -625 939 -613
rect 1351 613 1397 625
rect 1351 -613 1357 613
rect 1391 -613 1397 613
rect 1351 -625 1397 -613
rect 1809 613 1855 625
rect 1809 -613 1815 613
rect 1849 -613 1855 613
rect 1809 -625 1855 -613
rect 2267 613 2313 625
rect 2267 -613 2273 613
rect 2307 -613 2313 613
rect 2267 -625 2313 -613
rect 2725 613 2771 625
rect 2725 -613 2731 613
rect 2765 -613 2771 613
rect 2725 -625 2771 -613
rect 3183 613 3229 625
rect 3183 -613 3189 613
rect 3223 -613 3229 613
rect 3183 -625 3229 -613
rect 3641 613 3687 625
rect 3641 -613 3647 613
rect 3681 -613 3687 613
rect 3641 -625 3687 -613
rect -3631 -663 -3239 -657
rect -3631 -697 -3619 -663
rect -3251 -697 -3239 -663
rect -3631 -703 -3239 -697
rect -3173 -663 -2781 -657
rect -3173 -697 -3161 -663
rect -2793 -697 -2781 -663
rect -3173 -703 -2781 -697
rect -2715 -663 -2323 -657
rect -2715 -697 -2703 -663
rect -2335 -697 -2323 -663
rect -2715 -703 -2323 -697
rect -2257 -663 -1865 -657
rect -2257 -697 -2245 -663
rect -1877 -697 -1865 -663
rect -2257 -703 -1865 -697
rect -1799 -663 -1407 -657
rect -1799 -697 -1787 -663
rect -1419 -697 -1407 -663
rect -1799 -703 -1407 -697
rect -1341 -663 -949 -657
rect -1341 -697 -1329 -663
rect -961 -697 -949 -663
rect -1341 -703 -949 -697
rect -883 -663 -491 -657
rect -883 -697 -871 -663
rect -503 -697 -491 -663
rect -883 -703 -491 -697
rect -425 -663 -33 -657
rect -425 -697 -413 -663
rect -45 -697 -33 -663
rect -425 -703 -33 -697
rect 33 -663 425 -657
rect 33 -697 45 -663
rect 413 -697 425 -663
rect 33 -703 425 -697
rect 491 -663 883 -657
rect 491 -697 503 -663
rect 871 -697 883 -663
rect 491 -703 883 -697
rect 949 -663 1341 -657
rect 949 -697 961 -663
rect 1329 -697 1341 -663
rect 949 -703 1341 -697
rect 1407 -663 1799 -657
rect 1407 -697 1419 -663
rect 1787 -697 1799 -663
rect 1407 -703 1799 -697
rect 1865 -663 2257 -657
rect 1865 -697 1877 -663
rect 2245 -697 2257 -663
rect 1865 -703 2257 -697
rect 2323 -663 2715 -657
rect 2323 -697 2335 -663
rect 2703 -697 2715 -663
rect 2323 -703 2715 -697
rect 2781 -663 3173 -657
rect 2781 -697 2793 -663
rect 3161 -697 3173 -663
rect 2781 -703 3173 -697
rect 3239 -663 3631 -657
rect 3239 -697 3251 -663
rect 3619 -697 3631 -663
rect 3239 -703 3631 -697
<< properties >>
string FIXED_BBOX -3778 -782 3778 782
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 6.25 l 2.0 m 1 nf 16 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
