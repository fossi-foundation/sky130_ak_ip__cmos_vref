magic
tech sky130A
magscale 1 2
timestamp 1713056482
<< pwell >>
rect -235 -1442 235 1442
<< psubdiff >>
rect -199 1372 -103 1406
rect 103 1372 199 1406
rect -199 1310 -165 1372
rect 165 1310 199 1372
rect -199 -1372 -165 -1310
rect 165 -1372 199 -1310
rect -199 -1406 -103 -1372
rect 103 -1406 199 -1372
<< psubdiffcont >>
rect -103 1372 103 1406
rect -199 -1310 -165 1310
rect 165 -1310 199 1310
rect -103 -1406 103 -1372
<< xpolycontact >>
rect -69 844 69 1276
rect -69 -1276 69 -844
<< xpolyres >>
rect -69 -844 69 844
<< locali >>
rect -199 1372 -103 1406
rect 103 1372 199 1406
rect -199 1310 -165 1372
rect 165 1310 199 1372
rect -199 -1372 -165 -1310
rect 165 -1372 199 -1310
rect -199 -1406 -103 -1372
rect 103 -1406 199 -1372
<< viali >>
rect -53 861 53 1258
rect -53 -1258 53 -861
<< metal1 >>
rect -59 1258 59 1270
rect -59 861 -53 1258
rect 53 861 59 1258
rect -59 849 59 861
rect -59 -861 59 -849
rect -59 -1258 -53 -861
rect 53 -1258 59 -861
rect -59 -1270 59 -1258
<< properties >>
string FIXED_BBOX -182 -1389 182 1389
string gencell sky130_fd_pr__res_xhigh_po_0p69
string library sky130
string parameters w 0.690 l 8.6 m 1 nx 1 wmin 0.690 lmin 0.50 rho 2000 val 25.473k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.690 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
