magic
tech sky130A
magscale 1 2
timestamp 1713118989
use sky130_fd_pr__res_xhigh_po_0p69_2G52HS  sky130_fd_pr__res_xhigh_po_0p69_2G52HS_0
timestamp 1713051387
transform 1 0 4432 0 1 -813
box -352 -927 352 927
use sky130_fd_pr__res_xhigh_po_0p69_D5BT6X  sky130_fd_pr__res_xhigh_po_0p69_D5BT6X_0
timestamp 1713051387
transform 1 0 4654 0 1 -3133
box -1054 -927 1054 927
use sky130_fd_pr__res_xhigh_po_0p69_H5FMR6  sky130_fd_pr__res_xhigh_po_0p69_H5FMR6_0
timestamp 1713051387
transform 1 0 3835 0 1 -813
box -235 -927 235 927
use sky130_fd_pr__res_xhigh_po_0p69_H5TM75  sky130_fd_pr__res_xhigh_po_0p69_H5TM75_0
timestamp 1713051387
transform 1 0 5386 0 1 -813
box -586 -927 586 927
use sky130_fd_pr__nfet_01v8_J222PV  XM1
timestamp 1713050122
transform 1 0 2605 0 1 -1030
box -625 -710 625 710
use sky130_fd_pr__nfet_01v8_J222PV  XM2
timestamp 1713050122
transform 1 0 1345 0 1 -1030
box -625 -710 625 710
use sky130_fd_pr__nfet_01v8_J222PV  XM3
timestamp 1713050122
transform 1 0 1345 0 1 -2910
box -625 -710 625 710
use sky130_fd_pr__nfet_01v8_J222PV  XM4
timestamp 1713050122
transform 1 0 2605 0 1 -2910
box -625 -710 625 710
<< end >>
