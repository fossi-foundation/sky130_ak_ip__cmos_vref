magic
tech sky130A
timestamp 1713045697
<< pwell >>
rect -1406 -205 1406 205
<< nmos >>
rect -1308 -100 -808 100
rect -779 -100 -279 100
rect -250 -100 250 100
rect 279 -100 779 100
rect 808 -100 1308 100
<< ndiff >>
rect -1337 94 -1308 100
rect -1337 -94 -1331 94
rect -1314 -94 -1308 94
rect -1337 -100 -1308 -94
rect -808 94 -779 100
rect -808 -94 -802 94
rect -785 -94 -779 94
rect -808 -100 -779 -94
rect -279 94 -250 100
rect -279 -94 -273 94
rect -256 -94 -250 94
rect -279 -100 -250 -94
rect 250 94 279 100
rect 250 -94 256 94
rect 273 -94 279 94
rect 250 -100 279 -94
rect 779 94 808 100
rect 779 -94 785 94
rect 802 -94 808 94
rect 779 -100 808 -94
rect 1308 94 1337 100
rect 1308 -94 1314 94
rect 1331 -94 1337 94
rect 1308 -100 1337 -94
<< ndiffc >>
rect -1331 -94 -1314 94
rect -802 -94 -785 94
rect -273 -94 -256 94
rect 256 -94 273 94
rect 785 -94 802 94
rect 1314 -94 1331 94
<< psubdiff >>
rect -1388 170 -1340 187
rect 1340 170 1388 187
rect -1388 139 -1371 170
rect 1371 139 1388 170
rect -1388 -170 -1371 -139
rect 1371 -170 1388 -139
rect -1388 -187 -1340 -170
rect 1340 -187 1388 -170
<< psubdiffcont >>
rect -1340 170 1340 187
rect -1388 -139 -1371 139
rect 1371 -139 1388 139
rect -1340 -187 1340 -170
<< poly >>
rect -1308 136 -808 144
rect -1308 119 -1300 136
rect -816 119 -808 136
rect -1308 100 -808 119
rect -779 136 -279 144
rect -779 119 -771 136
rect -287 119 -279 136
rect -779 100 -279 119
rect -250 136 250 144
rect -250 119 -242 136
rect 242 119 250 136
rect -250 100 250 119
rect 279 136 779 144
rect 279 119 287 136
rect 771 119 779 136
rect 279 100 779 119
rect 808 136 1308 144
rect 808 119 816 136
rect 1300 119 1308 136
rect 808 100 1308 119
rect -1308 -119 -808 -100
rect -1308 -136 -1300 -119
rect -816 -136 -808 -119
rect -1308 -144 -808 -136
rect -779 -119 -279 -100
rect -779 -136 -771 -119
rect -287 -136 -279 -119
rect -779 -144 -279 -136
rect -250 -119 250 -100
rect -250 -136 -242 -119
rect 242 -136 250 -119
rect -250 -144 250 -136
rect 279 -119 779 -100
rect 279 -136 287 -119
rect 771 -136 779 -119
rect 279 -144 779 -136
rect 808 -119 1308 -100
rect 808 -136 816 -119
rect 1300 -136 1308 -119
rect 808 -144 1308 -136
<< polycont >>
rect -1300 119 -816 136
rect -771 119 -287 136
rect -242 119 242 136
rect 287 119 771 136
rect 816 119 1300 136
rect -1300 -136 -816 -119
rect -771 -136 -287 -119
rect -242 -136 242 -119
rect 287 -136 771 -119
rect 816 -136 1300 -119
<< locali >>
rect -1388 170 -1340 187
rect 1340 170 1388 187
rect -1388 139 -1371 170
rect 1371 139 1388 170
rect -1308 119 -1300 136
rect -816 119 -808 136
rect -779 119 -771 136
rect -287 119 -279 136
rect -250 119 -242 136
rect 242 119 250 136
rect 279 119 287 136
rect 771 119 779 136
rect 808 119 816 136
rect 1300 119 1308 136
rect -1331 94 -1314 102
rect -1331 -102 -1314 -94
rect -802 94 -785 102
rect -802 -102 -785 -94
rect -273 94 -256 102
rect -273 -102 -256 -94
rect 256 94 273 102
rect 256 -102 273 -94
rect 785 94 802 102
rect 785 -102 802 -94
rect 1314 94 1331 102
rect 1314 -102 1331 -94
rect -1308 -136 -1300 -119
rect -816 -136 -808 -119
rect -779 -136 -771 -119
rect -287 -136 -279 -119
rect -250 -136 -242 -119
rect 242 -136 250 -119
rect 279 -136 287 -119
rect 771 -136 779 -119
rect 808 -136 816 -119
rect 1300 -136 1308 -119
rect -1388 -170 -1371 -139
rect 1371 -170 1388 -139
rect -1388 -187 -1340 -170
rect 1340 -187 1388 -170
<< viali >>
rect -1300 119 -816 136
rect -771 119 -287 136
rect -242 119 242 136
rect 287 119 771 136
rect 816 119 1300 136
rect -1331 -94 -1314 94
rect -802 -94 -785 94
rect -273 -94 -256 94
rect 256 -94 273 94
rect 785 -94 802 94
rect 1314 -94 1331 94
rect -1300 -136 -816 -119
rect -771 -136 -287 -119
rect -242 -136 242 -119
rect 287 -136 771 -119
rect 816 -136 1300 -119
<< metal1 >>
rect -1306 136 -810 139
rect -1306 119 -1300 136
rect -816 119 -810 136
rect -1306 116 -810 119
rect -777 136 -281 139
rect -777 119 -771 136
rect -287 119 -281 136
rect -777 116 -281 119
rect -248 136 248 139
rect -248 119 -242 136
rect 242 119 248 136
rect -248 116 248 119
rect 281 136 777 139
rect 281 119 287 136
rect 771 119 777 136
rect 281 116 777 119
rect 810 136 1306 139
rect 810 119 816 136
rect 1300 119 1306 136
rect 810 116 1306 119
rect -1334 94 -1311 100
rect -1334 -94 -1331 94
rect -1314 -94 -1311 94
rect -1334 -100 -1311 -94
rect -805 94 -782 100
rect -805 -94 -802 94
rect -785 -94 -782 94
rect -805 -100 -782 -94
rect -276 94 -253 100
rect -276 -94 -273 94
rect -256 -94 -253 94
rect -276 -100 -253 -94
rect 253 94 276 100
rect 253 -94 256 94
rect 273 -94 276 94
rect 253 -100 276 -94
rect 782 94 805 100
rect 782 -94 785 94
rect 802 -94 805 94
rect 782 -100 805 -94
rect 1311 94 1334 100
rect 1311 -94 1314 94
rect 1331 -94 1334 94
rect 1311 -100 1334 -94
rect -1306 -119 -810 -116
rect -1306 -136 -1300 -119
rect -816 -136 -810 -119
rect -1306 -139 -810 -136
rect -777 -119 -281 -116
rect -777 -136 -771 -119
rect -287 -136 -281 -119
rect -777 -139 -281 -136
rect -248 -119 248 -116
rect -248 -136 -242 -119
rect 242 -136 248 -119
rect -248 -139 248 -136
rect 281 -119 777 -116
rect 281 -136 287 -119
rect 771 -136 777 -119
rect 281 -139 777 -136
rect 810 -119 1306 -116
rect 810 -136 816 -119
rect 1300 -136 1306 -119
rect 810 -139 1306 -136
<< properties >>
string FIXED_BBOX -1379 -178 1379 178
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2.0 l 5.0 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
