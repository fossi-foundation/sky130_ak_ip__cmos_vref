magic
tech sky130A
timestamp 1713045697
<< pwell >>
rect -1098 -230 1098 230
<< nmos >>
rect -1000 -125 1000 125
<< ndiff >>
rect -1029 119 -1000 125
rect -1029 -119 -1023 119
rect -1006 -119 -1000 119
rect -1029 -125 -1000 -119
rect 1000 119 1029 125
rect 1000 -119 1006 119
rect 1023 -119 1029 119
rect 1000 -125 1029 -119
<< ndiffc >>
rect -1023 -119 -1006 119
rect 1006 -119 1023 119
<< psubdiff >>
rect -1080 195 -1032 212
rect 1032 195 1080 212
rect -1080 164 -1063 195
rect 1063 164 1080 195
rect -1080 -195 -1063 -164
rect 1063 -195 1080 -164
rect -1080 -212 -1032 -195
rect 1032 -212 1080 -195
<< psubdiffcont >>
rect -1032 195 1032 212
rect -1080 -164 -1063 164
rect 1063 -164 1080 164
rect -1032 -212 1032 -195
<< poly >>
rect -1000 161 1000 169
rect -1000 144 -992 161
rect 992 144 1000 161
rect -1000 125 1000 144
rect -1000 -144 1000 -125
rect -1000 -161 -992 -144
rect 992 -161 1000 -144
rect -1000 -169 1000 -161
<< polycont >>
rect -992 144 992 161
rect -992 -161 992 -144
<< locali >>
rect -1080 195 -1032 212
rect 1032 195 1080 212
rect -1080 164 -1063 195
rect 1063 164 1080 195
rect -1000 144 -992 161
rect 992 144 1000 161
rect -1023 119 -1006 127
rect -1023 -127 -1006 -119
rect 1006 119 1023 127
rect 1006 -127 1023 -119
rect -1000 -161 -992 -144
rect 992 -161 1000 -144
rect -1080 -195 -1063 -164
rect 1063 -195 1080 -164
rect -1080 -212 -1032 -195
rect 1032 -212 1080 -195
<< viali >>
rect -992 144 992 161
rect -1023 -119 -1006 119
rect 1006 -119 1023 119
rect -992 -161 992 -144
<< metal1 >>
rect -998 161 998 164
rect -998 144 -992 161
rect 992 144 998 161
rect -998 141 998 144
rect -1026 119 -1003 125
rect -1026 -119 -1023 119
rect -1006 -119 -1003 119
rect -1026 -125 -1003 -119
rect 1003 119 1026 125
rect 1003 -119 1006 119
rect 1023 -119 1026 119
rect 1003 -125 1026 -119
rect -998 -144 998 -141
rect -998 -161 -992 -144
rect 992 -161 998 -144
rect -998 -164 998 -161
<< properties >>
string FIXED_BBOX -1071 -203 1071 203
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2.5 l 20.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
