magic
tech sky130A
magscale 1 2
timestamp 1713116496
<< error_s >>
rect 2500 -926 2506 -920
rect 2694 -926 2700 -920
rect 2494 -932 2500 -926
rect 2700 -932 2706 -926
rect 2494 -1126 2500 -1120
rect 2700 -1126 2706 -1120
rect 2500 -1132 2506 -1126
rect 2694 -1132 2700 -1126
rect 5660 -1240 5666 -1234
rect 5854 -1240 5860 -1234
rect 5654 -1246 5660 -1240
rect 5860 -1246 5866 -1240
rect 4660 -1272 4666 -1266
rect 4666 -1278 4672 -1272
rect 5654 -1440 5660 -1435
rect 5860 -1440 5866 -1435
rect 5660 -1446 5666 -1440
rect 5854 -1446 5860 -1440
<< metal1 >>
rect 3160 220 3360 460
rect 720 0 2938 200
rect 720 -260 1676 -60
rect 1020 -580 1220 -260
rect 1476 -540 1676 -260
rect 2280 -560 2480 0
rect 2738 -562 2938 0
rect 1246 -912 1446 -906
rect 1246 -1118 1446 -1112
rect 862 -1294 1092 -1276
rect 862 -1494 880 -1294
rect 1080 -1494 1092 -1294
rect 862 -1510 1092 -1494
rect 1638 -1294 1838 -1288
rect 1638 -1500 1838 -1494
rect 2118 -1302 2330 -1296
rect 2118 -1500 2124 -1302
rect 2324 -1500 2330 -1302
rect 2118 -1508 2330 -1500
rect 2890 -1302 3090 -1296
rect 2890 -1508 3090 -1500
rect 1640 -2420 1840 -2414
rect 2900 -2420 3100 -2414
rect 854 -2620 860 -2420
rect 1060 -2620 1066 -2420
rect 2094 -2620 2100 -2420
rect 2300 -2620 2306 -2420
rect 1640 -2626 1840 -2620
rect 2900 -2626 3100 -2620
rect 3160 -2499 3361 220
rect 3420 -1300 3620 460
rect 3736 -808 3936 -198
rect 4214 -390 4652 -190
rect 4942 -378 5342 -178
rect 5424 -372 5824 -172
rect 3736 -1008 4394 -808
rect 4194 -1278 4394 -1008
rect 4460 -1272 5120 -1260
rect 3720 -1300 3920 -1296
rect 3420 -1302 3920 -1300
rect 3420 -1500 3720 -1302
rect 4188 -1478 4194 -1278
rect 4394 -1478 4400 -1278
rect 4460 -1472 4466 -1272
rect 4666 -1460 5120 -1272
rect 5180 -1456 5580 -1256
rect 4666 -1472 4672 -1460
rect 4194 -1492 4394 -1478
rect 3720 -1508 3920 -1500
rect 5660 -2414 5860 -1440
rect 5660 -2420 5880 -2414
rect 5660 -2480 5680 -2420
rect 1240 -2700 1440 -2694
rect 3160 -2700 3920 -2499
rect 3980 -2680 4380 -2480
rect 4460 -2680 4860 -2480
rect 4920 -2680 5320 -2480
rect 5380 -2620 5680 -2480
rect 5380 -2626 5880 -2620
rect 5380 -2680 5860 -2626
rect 2494 -2900 2500 -2700
rect 2700 -2900 2706 -2700
rect 3154 -2900 3160 -2700
rect 3360 -2900 3366 -2700
rect 1240 -2906 1440 -2900
rect 1020 -3700 1220 -3400
rect 1460 -3700 1660 -3400
rect 720 -3900 1660 -3700
rect 2300 -3980 2500 -3420
rect 2760 -3980 2960 -3420
rect 3740 -3780 4140 -3580
rect 4220 -3760 4620 -3560
rect 4680 -3760 5080 -3560
rect 5160 -3760 5560 -3560
rect 720 -4180 2960 -3980
<< via1 >>
rect 1246 -1112 1446 -912
rect 2500 -1126 2700 -926
rect 880 -1494 1080 -1294
rect 1638 -1494 1838 -1294
rect 2124 -1500 2324 -1302
rect 2890 -1500 3090 -1302
rect 860 -2620 1060 -2420
rect 1640 -2620 1840 -2420
rect 2100 -2620 2300 -2420
rect 2900 -2620 3100 -2420
rect 3720 -1500 3920 -1302
rect 4194 -1478 4394 -1278
rect 4466 -1472 4666 -1272
rect 5660 -1440 5860 -1240
rect 5680 -2620 5880 -2420
rect 1240 -2900 1440 -2700
rect 2500 -2900 2700 -2700
rect 3160 -2900 3360 -2700
<< metal2 >>
rect 1240 -880 4660 -680
rect 1240 -912 1446 -880
rect 1240 -940 1246 -912
rect 1446 -1112 1452 -912
rect 1246 -1140 1440 -1112
rect 1640 -1126 2500 -926
rect 2700 -1126 4380 -926
rect 862 -1294 1092 -1276
rect 1640 -1294 1840 -1126
rect 4180 -1272 4380 -1126
rect 4460 -1272 4660 -880
rect 4180 -1278 4394 -1272
rect 862 -1494 880 -1294
rect 1080 -1494 1638 -1294
rect 1838 -1494 1844 -1294
rect 2118 -1302 2330 -1296
rect 862 -1510 1092 -1494
rect 1248 -1500 1448 -1494
rect 1640 -1500 1840 -1494
rect 2118 -1500 2124 -1302
rect 2324 -1500 2890 -1302
rect 3090 -1500 3720 -1302
rect 3920 -1500 3926 -1302
rect 4180 -1478 4194 -1278
rect 4180 -1480 4394 -1478
rect 4194 -1500 4394 -1480
rect 4460 -1472 4466 -1272
rect 4666 -1472 4680 -1320
rect 5656 -1435 5660 -1245
rect 5860 -1435 5864 -1245
rect 4460 -1640 4680 -1472
rect 4480 -1840 4680 -1640
rect 1320 -2040 4680 -1840
rect 1320 -2360 1520 -2040
rect 860 -2420 1060 -2414
rect 1300 -2420 1520 -2360
rect 2100 -2420 2300 -2414
rect 1060 -2620 1640 -2420
rect 1840 -2620 1846 -2420
rect 2300 -2620 2900 -2420
rect 3100 -2620 5680 -2420
rect 5880 -2620 5886 -2420
rect 860 -2626 1060 -2620
rect 2100 -2626 2320 -2620
rect 2120 -2700 2320 -2626
rect 1220 -2900 1240 -2700
rect 1440 -2900 2320 -2700
rect 2500 -2700 2700 -2694
rect 3160 -2700 3360 -2694
rect 2700 -2900 3160 -2700
rect 3360 -2900 3380 -2700
rect 2500 -2906 2700 -2900
rect 3160 -2906 3360 -2900
use sky130_fd_pr__res_xhigh_po_0p69_2G52HS  sky130_fd_pr__res_xhigh_po_0p69_2G52HS_0
timestamp 1713051387
transform 1 0 4432 0 1 -813
box -352 -927 352 927
use sky130_fd_pr__res_xhigh_po_0p69_D5BT6X  sky130_fd_pr__res_xhigh_po_0p69_D5BT6X_0
timestamp 1713051387
transform 1 0 4654 0 1 -3133
box -1054 -927 1054 927
use sky130_fd_pr__res_xhigh_po_0p69_H5FMR6  sky130_fd_pr__res_xhigh_po_0p69_H5FMR6_0
timestamp 1713051387
transform 1 0 3835 0 1 -813
box -235 -927 235 927
use sky130_fd_pr__res_xhigh_po_0p69_H5TM75  sky130_fd_pr__res_xhigh_po_0p69_H5TM75_0
timestamp 1713051387
transform 1 0 5386 0 1 -813
box -586 -927 586 927
use sky130_fd_pr__nfet_01v8_J222PV  XM1
timestamp 1713050122
transform 1 0 2605 0 1 -1030
box -625 -710 625 710
use sky130_fd_pr__nfet_01v8_J222PV  XM2
timestamp 1713050122
transform 1 0 1345 0 1 -1030
box -625 -710 625 710
use sky130_fd_pr__nfet_01v8_J222PV  XM3
timestamp 1713050122
transform 1 0 1345 0 1 -2910
box -625 -710 625 710
use sky130_fd_pr__nfet_01v8_J222PV  XM4
timestamp 1713050122
transform 1 0 2605 0 1 -2910
box -625 -710 625 710
<< labels >>
flabel metal1 720 -260 920 -60 0 FreeSans 256 0 0 0 trim1
port 5 nsew
flabel metal1 720 -3900 920 -3700 0 FreeSans 256 0 0 0 trim2
port 3 nsew
flabel metal1 720 -4180 920 -3980 0 FreeSans 256 0 0 0 trim3
port 4 nsew
flabel metal1 3420 260 3620 460 0 FreeSans 256 0 0 0 A
port 1 nsew
flabel metal1 3160 260 3360 460 0 FreeSans 256 0 0 0 B
port 6 nsew
flabel metal1 720 0 920 200 0 FreeSans 256 0 0 0 trim0
port 2 nsew
<< end >>
