magic
tech sky130A
magscale 1 2
timestamp 1716165657
<< metal1 >>
rect 5700 4800 11200 5000
rect 5700 4619 5900 4800
rect 6000 4706 10892 4770
rect 8200 4619 8400 4706
rect 11000 4619 11200 4800
rect 5700 3619 5944 4619
rect 8048 3619 8400 4619
rect 5700 3500 5900 3619
rect 8200 3532 8400 3619
rect 6000 3468 8400 3532
rect 8200 3400 8400 3468
rect 5700 3360 8400 3400
rect 5700 3240 8240 3360
rect 8360 3240 8400 3360
rect 5700 3200 8400 3240
rect 8500 3619 8844 4619
rect 10948 3619 11200 4619
rect 8500 3391 8700 3619
rect 8900 3468 10892 3532
rect 8500 3200 8844 3391
rect 8900 3360 9060 3468
rect 8900 3240 8920 3360
rect 9040 3240 9060 3360
rect 8900 3220 9060 3240
rect 11000 3220 11200 3619
rect 6000 3146 7992 3152
rect 6000 3094 6006 3146
rect 7986 3094 7992 3146
rect 6000 3088 7992 3094
rect 5880 3005 5944 3010
rect 5880 1017 5886 3005
rect 5938 1017 5944 3005
rect 5880 1010 5944 1017
rect 8048 1240 8176 3200
rect 8280 3140 8520 3160
rect 8280 2940 8300 3140
rect 8500 2940 8520 3140
rect 8280 2920 8520 2940
rect 8048 1220 8260 1240
rect 8048 1020 8120 1220
rect 8048 1010 8260 1020
rect 8120 1000 8260 1010
rect 6000 900 7992 932
rect 8300 900 8500 2920
rect 8716 1240 8844 3200
rect 8900 3146 10892 3152
rect 8900 3094 8906 3146
rect 10886 3094 10892 3146
rect 8900 3088 10892 3094
rect 8540 1220 8844 1240
rect 8540 1020 8560 1220
rect 8700 1020 8844 1220
rect 8540 1010 8844 1020
rect 10948 3004 11012 3010
rect 10948 1016 10954 3004
rect 11006 1016 11012 3004
rect 10948 1010 11012 1016
rect 8540 1000 8720 1010
rect 8900 900 10892 932
rect 5700 700 10900 900
rect 8098 660 8341 661
rect 8098 641 9660 660
rect 8098 521 8119 641
rect 8319 540 9660 641
rect 8319 521 8341 540
rect 8098 501 8341 521
rect 8520 480 8760 500
rect 8520 460 8540 480
rect 5868 360 8540 460
rect 5868 -3400 5932 360
rect 8520 340 8540 360
rect 8740 340 8760 480
rect 8520 330 8760 340
rect 8520 320 9312 330
rect 8588 266 9312 320
rect 6010 257 8510 263
rect 6010 205 6016 257
rect 8394 205 8510 257
rect 6010 199 8510 205
rect 6010 -201 8510 -195
rect 6010 -253 6126 -201
rect 8504 -253 8510 -201
rect 6010 -259 8510 -253
rect 6010 -659 8510 -653
rect 6010 -711 6016 -659
rect 8394 -711 8510 -659
rect 6010 -717 8510 -711
rect 8588 -890 8716 266
rect 8855 182 8919 188
rect 8855 -806 8861 182
rect 8913 -806 8919 182
rect 8855 -812 8919 -806
rect 9368 182 9432 188
rect 9368 -806 9374 182
rect 9426 -806 9432 182
rect 9368 -812 9432 -806
rect 9540 -824 9660 540
rect 11040 -680 11200 3220
rect 10920 -700 11200 -680
rect 8588 -954 9312 -890
rect 9540 -952 10710 -824
rect 10920 -940 10940 -700
rect 11180 -940 11200 -700
rect 6010 -1117 8510 -1111
rect 6010 -1169 6126 -1117
rect 8504 -1169 8510 -1117
rect 6010 -1175 8510 -1169
rect 6010 -1575 8510 -1569
rect 6010 -1627 6016 -1575
rect 8394 -1627 8510 -1575
rect 6010 -1633 8510 -1627
rect 6010 -2033 8510 -2027
rect 6010 -2085 6126 -2033
rect 8504 -2085 8510 -2033
rect 6010 -2091 8510 -2085
rect 8588 -2260 8716 -954
rect 10920 -960 11200 -940
rect 9280 -1080 9520 -1060
rect 9280 -1280 9300 -1080
rect 9500 -1280 9520 -1080
rect 9280 -1300 9520 -1280
rect 9300 -2200 9500 -1300
rect 9568 -1898 9632 -1008
rect 9568 -2154 9574 -1898
rect 9626 -2154 9632 -1898
rect 10787 -1020 10915 -1008
rect 10787 -1040 11200 -1020
rect 10787 -1280 10940 -1040
rect 11180 -1280 11200 -1040
rect 10787 -1300 11200 -1280
rect 10787 -1898 10915 -1300
rect 9568 -2160 9632 -2154
rect 9710 -2200 10710 -2056
rect 8588 -2280 8940 -2260
rect 8588 -2480 8720 -2280
rect 8920 -2480 8940 -2280
rect 6010 -2491 8510 -2485
rect 6010 -2543 6016 -2491
rect 8394 -2543 8510 -2491
rect 6010 -2549 8510 -2543
rect 8588 -2500 8940 -2480
rect 9300 -2300 10710 -2200
rect 10787 -2154 10794 -1898
rect 10846 -2154 10915 -1898
rect 9300 -2490 9500 -2300
rect 9700 -2354 10692 -2348
rect 9700 -2406 9706 -2354
rect 10686 -2406 10692 -2354
rect 9700 -2412 10692 -2406
rect 10787 -2490 10915 -2154
rect 6010 -2949 8510 -2943
rect 6010 -3001 6126 -2949
rect 8504 -3001 8510 -2949
rect 6010 -3007 8510 -3001
rect 8588 -3400 8716 -2500
rect 6010 -3407 8510 -3401
rect 6010 -3459 6016 -3407
rect 8394 -3459 8510 -3407
rect 6010 -3465 8510 -3459
rect 9300 -3490 9644 -2490
rect 10748 -3490 10915 -2490
rect 8300 -3520 8900 -3500
rect 8300 -3580 8320 -3520
rect 8680 -3580 8900 -3520
rect 8300 -3600 8900 -3580
rect 8700 -3700 8900 -3600
rect 9300 -3700 9500 -3490
rect 9700 -3574 10692 -3568
rect 9700 -3626 9706 -3574
rect 10686 -3626 10692 -3574
rect 9700 -3632 10692 -3626
<< via1 >>
rect 8240 3240 8360 3360
rect 8920 3240 9040 3360
rect 6006 3094 7986 3146
rect 5886 1017 5938 3005
rect 8300 2940 8500 3140
rect 8120 1020 8260 1220
rect 8906 3094 10886 3146
rect 8560 1020 8700 1220
rect 10954 1016 11006 3004
rect 8119 521 8319 641
rect 8540 340 8740 480
rect 6016 205 8394 257
rect 6126 -253 8504 -201
rect 6016 -711 8394 -659
rect 8861 -806 8913 182
rect 9374 -806 9426 182
rect 10940 -940 11180 -700
rect 6126 -1169 8504 -1117
rect 6016 -1627 8394 -1575
rect 6126 -2085 8504 -2033
rect 9300 -1280 9500 -1080
rect 9574 -2154 9626 -1898
rect 10940 -1280 11180 -1040
rect 8720 -2480 8920 -2280
rect 6016 -2543 8394 -2491
rect 10794 -2154 10846 -1898
rect 9706 -2406 10686 -2354
rect 6126 -3001 8504 -2949
rect 6016 -3459 8394 -3407
rect 8320 -3580 8680 -3520
rect 9706 -3626 10686 -3574
<< metal2 >>
rect 8220 3360 8380 3380
rect 8900 3360 9060 3380
rect 8220 3240 8240 3360
rect 8360 3240 8920 3360
rect 9040 3240 9060 3360
rect 8220 3220 8380 3240
rect 8900 3220 9060 3240
rect 8280 3152 8520 3160
rect 6000 3146 10892 3152
rect 6000 3094 6006 3146
rect 7986 3140 8906 3146
rect 7986 3094 8300 3140
rect 6000 3088 8300 3094
rect 5816 3005 5944 3010
rect 5816 1017 5886 3005
rect 5938 1017 5944 3005
rect 8280 2940 8300 3088
rect 8500 3094 8906 3140
rect 10886 3094 10892 3146
rect 8500 3088 10892 3094
rect 8500 2940 8520 3088
rect 8280 2920 8520 2940
rect 10948 3004 11076 3010
rect 5816 664 5944 1017
rect 8120 1220 8260 1240
rect 5816 536 6010 664
rect 8120 661 8260 1020
rect 8540 1220 8720 1240
rect 8540 1020 8560 1220
rect 8700 1020 8720 1220
rect 8540 1000 8720 1020
rect 10948 1016 10954 3004
rect 11006 1016 11076 3004
rect 5882 263 6010 536
rect 8098 641 8341 661
rect 8098 521 8119 641
rect 8319 521 8341 641
rect 8098 501 8341 521
rect 8560 500 8700 1000
rect 10948 664 11076 1016
rect 9376 536 11076 664
rect 8520 480 8760 500
rect 8520 340 8540 480
rect 8740 340 8760 480
rect 8520 320 8760 340
rect 5882 257 8400 263
rect 5882 205 6016 257
rect 8394 205 8400 257
rect 5882 199 8400 205
rect 5882 -653 6010 199
rect 9376 188 9504 536
rect 8791 182 8919 188
rect 6120 -201 8638 -195
rect 6120 -253 6126 -201
rect 8504 -253 8638 -201
rect 6120 -259 8638 -253
rect 5882 -659 8400 -653
rect 5882 -711 6016 -659
rect 8394 -711 8400 -659
rect 5882 -717 8400 -711
rect 5882 -1569 6010 -717
rect 8510 -1111 8638 -259
rect 6120 -1117 8638 -1111
rect 6120 -1169 6126 -1117
rect 8504 -1169 8638 -1117
rect 6120 -1175 8638 -1169
rect 5882 -1575 8400 -1569
rect 5882 -1627 6016 -1575
rect 8394 -1627 8400 -1575
rect 5882 -1633 8400 -1627
rect 5882 -2485 6010 -1633
rect 8510 -2026 8638 -1175
rect 8791 -806 8861 182
rect 8913 -806 8919 182
rect 8791 -1060 8919 -806
rect 9368 182 9504 188
rect 9368 -806 9374 182
rect 9426 -806 9504 182
rect 9368 -811 9504 -806
rect 10920 -700 11200 -680
rect 10920 -940 10940 -700
rect 11180 -940 11200 -700
rect 10920 -960 11200 -940
rect 10920 -1040 11200 -1020
rect 8791 -1080 9520 -1060
rect 8791 -1280 9300 -1080
rect 9500 -1280 9520 -1080
rect 8791 -1300 9520 -1280
rect 10920 -1280 10940 -1040
rect 11180 -1280 11200 -1040
rect 10920 -1300 11200 -1280
rect 6120 -2033 8638 -2026
rect 6120 -2085 6126 -2033
rect 8504 -2085 8638 -2033
rect 6120 -2090 8638 -2085
rect 5882 -2491 8400 -2485
rect 5882 -2543 6016 -2491
rect 8394 -2543 8400 -2491
rect 5882 -2549 8400 -2543
rect 5882 -3401 6010 -2549
rect 8510 -2943 8638 -2090
rect 9568 -1898 9632 -1892
rect 9568 -2154 9574 -1898
rect 9626 -2096 9632 -1898
rect 10788 -1898 10852 -1892
rect 10788 -2096 10794 -1898
rect 9626 -2154 10794 -2096
rect 10846 -2154 10852 -1898
rect 9568 -2160 10852 -2154
rect 8700 -2280 8940 -2260
rect 8700 -2480 8720 -2280
rect 8920 -2348 8940 -2280
rect 8920 -2354 10945 -2348
rect 8920 -2406 9706 -2354
rect 10686 -2406 10945 -2354
rect 8920 -2412 10945 -2406
rect 8920 -2480 8940 -2412
rect 8700 -2500 8940 -2480
rect 6120 -2949 8638 -2943
rect 6120 -3001 6126 -2949
rect 8504 -3001 8638 -2949
rect 6120 -3007 8638 -3001
rect 5882 -3407 8400 -3401
rect 5882 -3459 6016 -3407
rect 8394 -3459 8400 -3407
rect 5882 -3465 8400 -3459
rect 8510 -3500 8638 -3007
rect 8300 -3520 8700 -3500
rect 8300 -3580 8320 -3520
rect 8680 -3580 8700 -3520
rect 10881 -3568 10945 -2412
rect 8300 -3600 8700 -3580
rect 9700 -3574 10945 -3568
rect 9700 -3626 9706 -3574
rect 10686 -3626 10945 -3574
rect 9700 -3632 10945 -3626
<< via2 >>
rect 10940 -940 11180 -700
rect 10940 -1280 11180 -1040
<< metal3 >>
rect 10920 -700 11200 -680
rect 10920 -940 10940 -700
rect 11180 -940 11200 -700
rect 10920 -960 11200 -940
rect 10920 -1040 11200 -1020
rect 10920 -1280 10940 -1040
rect 11180 -1280 11200 -1040
rect 10920 -1300 11200 -1280
<< via3 >>
rect 10940 -940 11180 -700
rect 10940 -1280 11180 -1040
<< metal4 >>
rect 9740 -560 10739 442
rect 10200 -660 10300 -560
rect 10200 -760 10810 -660
rect 10972 -680 11068 -588
rect 10710 -1100 10810 -760
rect 10920 -700 11200 -680
rect 10920 -940 10940 -700
rect 11180 -940 11200 -700
rect 10920 -960 11200 -940
rect 10920 -1040 11200 -1020
rect 10920 -1100 10940 -1040
rect 10710 -1200 10940 -1100
rect 10920 -1280 10940 -1200
rect 11180 -1280 11200 -1040
rect 10920 -1300 11200 -1280
use sky130_fd_pr__nfet_01v8_QTPFY2  sky130_fd_pr__nfet_01v8_QTPFY2_0
timestamp 1713212409
transform 0 1 7260 -1 0 -1601
box -1999 -1460 1999 1460
use sky130_fd_pr__cap_mim_m3_1_VCAG9S  XC1
timestamp 1713045697
transform 1 0 10386 0 1 -60
box -686 -540 686 540
use sky130_fd_pr__nfet_01v8_QGRVRG  XM4
timestamp 1713045697
transform 1 0 9116 0 1 -312
box -396 -710 396 710
use sky130_fd_pr__nfet_01v8_ME6MQD  XM5
timestamp 1713045697
transform 1 0 6996 0 1 2010
box -1196 -1210 1196 1210
use sky130_fd_pr__nfet_01v8_ME6MQD  XM6
timestamp 1713045697
transform 1 0 9896 0 1 2010
box -1196 -1210 1196 1210
use sky130_fd_pr__pfet_01v8_6H4ZLK  XM7
timestamp 1716081177
transform 1 0 6996 0 1 4119
box -1196 -719 1196 719
use sky130_fd_pr__pfet_01v8_6H4ZLK  XM8
timestamp 1716081177
transform 1 0 9896 0 1 4119
box -1196 -719 1196 719
use sky130_fd_pr__nfet_01v8_TTEWAE  XM10
timestamp 1713212409
transform 0 -1 10210 1 0 -1504
box -696 -710 696 710
use sky130_fd_pr__nfet_01v8_BSH2JQ  XM11
timestamp 1713212409
transform -1 0 10196 0 -1 -2990
box -696 -710 696 710
<< labels >>
flabel metal1 5700 3500 5900 3700 0 FreeSans 256 0 0 0 vdd
port 0 nsew
flabel metal1 5700 3200 5900 3400 0 FreeSans 256 0 0 0 pbias
port 1 nsew
flabel metal1 5700 700 5900 900 0 FreeSans 256 0 0 0 nbias
port 2 nsew
flabel metal1 8700 -3700 8900 -3500 0 FreeSans 256 0 0 0 vx
port 3 nsew
flabel metal1 9300 -3700 9500 -3500 0 FreeSans 256 0 0 0 vss
port 4 nsew
<< end >>
