magic
tech sky130A
magscale 1 2
timestamp 1713045697
<< nwell >>
rect -1196 -5219 1196 5219
<< pmos >>
rect -1000 -5000 1000 5000
<< pdiff >>
rect -1058 4988 -1000 5000
rect -1058 -4988 -1046 4988
rect -1012 -4988 -1000 4988
rect -1058 -5000 -1000 -4988
rect 1000 4988 1058 5000
rect 1000 -4988 1012 4988
rect 1046 -4988 1058 4988
rect 1000 -5000 1058 -4988
<< pdiffc >>
rect -1046 -4988 -1012 4988
rect 1012 -4988 1046 4988
<< nsubdiff >>
rect -1160 5149 -1064 5183
rect 1064 5149 1160 5183
rect -1160 5087 -1126 5149
rect 1126 5087 1160 5149
rect -1160 -5149 -1126 -5087
rect 1126 -5149 1160 -5087
rect -1160 -5183 -1064 -5149
rect 1064 -5183 1160 -5149
<< nsubdiffcont >>
rect -1064 5149 1064 5183
rect -1160 -5087 -1126 5087
rect 1126 -5087 1160 5087
rect -1064 -5183 1064 -5149
<< poly >>
rect -1000 5081 1000 5097
rect -1000 5047 -984 5081
rect 984 5047 1000 5081
rect -1000 5000 1000 5047
rect -1000 -5047 1000 -5000
rect -1000 -5081 -984 -5047
rect 984 -5081 1000 -5047
rect -1000 -5097 1000 -5081
<< polycont >>
rect -984 5047 984 5081
rect -984 -5081 984 -5047
<< locali >>
rect -1160 5149 -1064 5183
rect 1064 5149 1160 5183
rect -1160 5087 -1126 5149
rect 1126 5087 1160 5149
rect -1000 5047 -984 5081
rect 984 5047 1000 5081
rect -1046 4988 -1012 5004
rect -1046 -5004 -1012 -4988
rect 1012 4988 1046 5004
rect 1012 -5004 1046 -4988
rect -1000 -5081 -984 -5047
rect 984 -5081 1000 -5047
rect -1160 -5149 -1126 -5087
rect 1126 -5149 1160 -5087
rect -1160 -5183 -1064 -5149
rect 1064 -5183 1160 -5149
<< viali >>
rect -984 5047 984 5081
rect -1046 -4988 -1012 4988
rect 1012 -4988 1046 4988
rect -984 -5081 984 -5047
<< metal1 >>
rect -996 5081 996 5087
rect -996 5047 -984 5081
rect 984 5047 996 5081
rect -996 5041 996 5047
rect -1052 4988 -1006 5000
rect -1052 -4988 -1046 4988
rect -1012 -4988 -1006 4988
rect -1052 -5000 -1006 -4988
rect 1006 4988 1052 5000
rect 1006 -4988 1012 4988
rect 1046 -4988 1052 4988
rect 1006 -5000 1052 -4988
rect -996 -5047 996 -5041
rect -996 -5081 -984 -5047
rect 984 -5081 996 -5047
rect -996 -5087 996 -5081
<< properties >>
string FIXED_BBOX -1143 -5166 1143 5166
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 50.0 l 10.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
