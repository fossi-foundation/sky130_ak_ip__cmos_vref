magic
tech sky130A
magscale 1 2
timestamp 1713045697
<< error_p >>
rect -414 1186 -264 1228
rect 264 1186 414 1228
rect -414 1174 -246 1186
rect -212 1174 212 1186
rect 246 1174 414 1186
rect -360 1152 -175 1174
rect 175 1152 414 1174
rect -360 1140 414 1152
rect -360 1090 -272 1140
rect -222 1106 -212 1110
rect 184 1106 222 1110
rect -372 1078 -272 1090
rect -360 -1078 -348 1078
rect -326 -1078 -314 1078
rect -234 1004 -206 1106
rect 184 1082 234 1106
rect 326 1090 414 1140
rect -194 1078 234 1082
rect 314 1078 414 1090
rect -196 1072 234 1078
rect -200 1038 -174 1072
rect 174 1038 234 1072
rect -196 1032 196 1038
rect -194 1028 194 1032
rect 206 1004 234 1038
rect -222 1000 -212 1004
rect 212 1000 222 1004
rect -222 -1004 -212 -1000
rect 184 -1004 222 -1000
rect -360 -1086 -272 -1078
rect -360 -1128 -264 -1086
rect -234 -1106 -206 -1004
rect 184 -1028 234 -1004
rect -194 -1032 234 -1028
rect -196 -1038 234 -1032
rect -200 -1072 -174 -1038
rect 174 -1072 234 -1038
rect -196 -1078 196 -1072
rect -194 -1082 194 -1078
rect 206 -1106 234 -1072
rect 326 -1078 338 1078
rect 360 -1078 372 1078
rect 326 -1086 414 -1078
rect -222 -1110 -212 -1106
rect 212 -1110 222 -1106
rect 264 -1128 414 -1086
rect -360 -1140 -246 -1128
rect -212 -1140 212 -1128
rect 246 -1140 414 -1128
rect -360 -1162 -175 -1140
rect 175 -1162 414 -1140
rect -360 -1174 414 -1162
<< pwell >>
rect -1312 -2210 1312 2210
<< nmos >>
rect -1116 -2000 -716 2000
rect -658 1174 -258 2000
rect -200 1174 200 2000
rect 258 1174 658 2000
rect -658 -1174 -360 1174
rect -326 -1140 -258 1140
rect -200 1072 200 1140
rect -200 1038 -184 1072
rect 184 1038 200 1072
rect -200 -1038 200 1038
rect -200 -1072 -184 -1038
rect 184 -1072 200 -1038
rect -200 -1140 200 -1072
rect 258 -1140 326 1140
rect 360 -1174 658 1174
rect -658 -2000 -258 -1174
rect -200 -2000 200 -1174
rect 258 -2000 658 -1174
rect 716 -2000 1116 2000
<< ndiff >>
rect -1174 1988 -1116 2000
rect -1174 -1988 -1162 1988
rect -1128 -1988 -1116 1988
rect -1174 -2000 -1116 -1988
rect -716 1988 -658 2000
rect -716 -1988 -704 1988
rect -670 -1988 -658 1988
rect -258 1988 -200 2000
rect -258 1174 -246 1988
rect -212 1174 -200 1988
rect 200 1988 258 2000
rect 200 1174 212 1988
rect 246 1174 258 1988
rect 658 1988 716 2000
rect -258 -1140 -246 1140
rect -212 -1140 -200 1140
rect 200 -1140 212 1140
rect 246 -1140 258 1140
rect -716 -2000 -658 -1988
rect -258 -1988 -246 -1174
rect -212 -1988 -200 -1174
rect -258 -2000 -200 -1988
rect 200 -1988 212 -1174
rect 246 -1988 258 -1174
rect 200 -2000 258 -1988
rect 658 -1988 670 1988
rect 704 -1988 716 1988
rect 658 -2000 716 -1988
rect 1116 1988 1174 2000
rect 1116 -1988 1128 1988
rect 1162 -1988 1174 1988
rect 1116 -2000 1174 -1988
<< ndiffc >>
rect -1162 -1988 -1128 1988
rect -704 -1988 -670 1988
rect -246 1174 -212 1988
rect 212 1174 246 1988
rect -246 -1140 -212 1140
rect 212 -1140 246 1140
rect -246 -1988 -212 -1174
rect 212 -1988 246 -1174
rect 670 -1988 704 1988
rect 1128 -1988 1162 1988
<< psubdiff >>
rect -1276 2140 -1180 2174
rect 1180 2140 1276 2174
rect -1276 2078 -1242 2140
rect 1242 2078 1276 2140
rect -360 1140 -264 1174
rect 264 1140 360 1174
rect -360 1078 -326 1140
rect -360 -1140 -326 -1078
rect 326 1078 360 1140
rect 326 -1140 360 -1078
rect -360 -1174 -264 -1140
rect 264 -1174 360 -1140
rect -1276 -2140 -1242 -2078
rect 1242 -2140 1276 -2078
rect -1276 -2174 -1180 -2140
rect 1180 -2174 1276 -2140
<< psubdiffcont >>
rect -1180 2140 1180 2174
rect -1276 -2078 -1242 2078
rect -264 1140 264 1174
rect -360 -1078 -326 1078
rect 326 -1078 360 1078
rect -264 -1174 264 -1140
rect 1242 -2078 1276 2078
rect -1180 -2174 1180 -2140
<< poly >>
rect -1116 2072 -716 2088
rect -1116 2038 -1100 2072
rect -732 2038 -716 2072
rect -1116 2000 -716 2038
rect -658 2072 -258 2088
rect -658 2038 -642 2072
rect -274 2038 -258 2072
rect -658 2000 -258 2038
rect -200 2072 200 2088
rect -200 2038 -184 2072
rect 184 2038 200 2072
rect -200 2000 200 2038
rect 258 2072 658 2088
rect 258 2038 274 2072
rect 642 2038 658 2072
rect 258 2000 658 2038
rect 716 2072 1116 2088
rect 716 2038 732 2072
rect 1100 2038 1116 2072
rect 716 2000 1116 2038
rect -1116 -2038 -716 -2000
rect -1116 -2072 -1100 -2038
rect -732 -2072 -716 -2038
rect -1116 -2088 -716 -2072
rect -658 -2038 -258 -2000
rect -658 -2072 -642 -2038
rect -274 -2072 -258 -2038
rect -658 -2088 -258 -2072
rect -200 -2038 200 -2000
rect -200 -2072 -184 -2038
rect 184 -2072 200 -2038
rect -200 -2088 200 -2072
rect 258 -2038 658 -2000
rect 258 -2072 274 -2038
rect 642 -2072 658 -2038
rect 258 -2088 658 -2072
rect 716 -2038 1116 -2000
rect 716 -2072 732 -2038
rect 1100 -2072 1116 -2038
rect 716 -2088 1116 -2072
<< polycont >>
rect -1100 2038 -732 2072
rect -642 2038 -274 2072
rect -184 2038 184 2072
rect 274 2038 642 2072
rect 732 2038 1100 2072
rect -184 1038 184 1072
rect -184 -1072 184 -1038
rect -1100 -2072 -732 -2038
rect -642 -2072 -274 -2038
rect -184 -2072 184 -2038
rect 274 -2072 642 -2038
rect 732 -2072 1100 -2038
<< locali >>
rect -1276 2140 -1180 2174
rect 1180 2140 1276 2174
rect -1276 2078 -1242 2140
rect 1242 2078 1276 2140
rect -1116 2038 -1100 2072
rect -732 2038 -716 2072
rect -658 2038 -642 2072
rect -274 2038 -258 2072
rect -200 2038 -184 2072
rect 184 2038 200 2072
rect 258 2038 274 2072
rect 642 2038 658 2072
rect 716 2038 732 2072
rect 1100 2038 1116 2072
rect -1162 1988 -1128 2004
rect -1162 -2004 -1128 -1988
rect -704 1988 -670 2004
rect -246 1988 -212 2004
rect 212 1988 246 2004
rect 670 1988 704 2004
rect -360 1140 -264 1174
rect 264 1140 360 1174
rect -360 1078 -326 1140
rect -360 -1140 -326 -1078
rect -200 1038 -184 1072
rect 184 1038 200 1072
rect -200 -1072 -184 -1038
rect 184 -1072 200 -1038
rect 326 1078 360 1140
rect 326 -1140 360 -1078
rect -360 -1174 -264 -1140
rect 264 -1174 360 -1140
rect -704 -2004 -670 -1988
rect -246 -2004 -212 -1988
rect 212 -2004 246 -1988
rect 670 -2004 704 -1988
rect 1128 1988 1162 2004
rect 1128 -2004 1162 -1988
rect -1116 -2072 -1100 -2038
rect -732 -2072 -716 -2038
rect -658 -2072 -642 -2038
rect -274 -2072 -258 -2038
rect -200 -2072 -184 -2038
rect 184 -2072 200 -2038
rect 258 -2072 274 -2038
rect 642 -2072 658 -2038
rect 716 -2072 732 -2038
rect 1100 -2072 1116 -2038
rect -1276 -2140 -1242 -2078
rect 1242 -2140 1276 -2078
rect -1276 -2174 -1180 -2140
rect 1180 -2174 1276 -2140
<< viali >>
rect -1100 2038 -732 2072
rect -642 2038 -274 2072
rect -184 2038 184 2072
rect 274 2038 642 2072
rect 732 2038 1100 2072
rect -1162 -1988 -1128 1988
rect -704 -1988 -670 1988
rect -246 1174 -212 1988
rect 212 1174 246 1988
rect -246 1140 -212 1174
rect 212 1140 246 1174
rect -246 -1140 -212 1140
rect -184 1038 184 1072
rect -184 -1072 184 -1038
rect 212 -1140 246 1140
rect -246 -1174 -212 -1140
rect 212 -1174 246 -1140
rect -246 -1988 -212 -1174
rect 212 -1988 246 -1174
rect 670 -1988 704 1988
rect 1128 -1988 1162 1988
rect -1100 -2072 -732 -2038
rect -642 -2072 -274 -2038
rect -184 -2072 184 -2038
rect 274 -2072 642 -2038
rect 732 -2072 1100 -2038
<< metal1 >>
rect -1112 2072 -720 2078
rect -1112 2038 -1100 2072
rect -732 2038 -720 2072
rect -1112 2032 -720 2038
rect -654 2072 -262 2078
rect -654 2038 -642 2072
rect -274 2038 -262 2072
rect -654 2032 -262 2038
rect -196 2072 196 2078
rect -196 2038 -184 2072
rect 184 2038 196 2072
rect -196 2032 196 2038
rect 262 2072 654 2078
rect 262 2038 274 2072
rect 642 2038 654 2072
rect 262 2032 654 2038
rect 720 2072 1112 2078
rect 720 2038 732 2072
rect 1100 2038 1112 2072
rect 720 2032 1112 2038
rect -1168 1988 -1122 2000
rect -1168 -1988 -1162 1988
rect -1128 -1988 -1122 1988
rect -1168 -2000 -1122 -1988
rect -710 1988 -664 2000
rect -710 -1988 -704 1988
rect -670 -1988 -664 1988
rect -710 -2000 -664 -1988
rect -252 1988 -206 2000
rect -252 -1988 -246 1988
rect -212 -1988 -206 1988
rect 206 1988 252 2000
rect -196 1072 196 1078
rect -196 1038 -184 1072
rect 184 1038 196 1072
rect -196 1032 196 1038
rect -196 -1038 196 -1032
rect -196 -1072 -184 -1038
rect 184 -1072 196 -1038
rect -196 -1078 196 -1072
rect -252 -2000 -206 -1988
rect 206 -1988 212 1988
rect 246 -1988 252 1988
rect 206 -2000 252 -1988
rect 664 1988 710 2000
rect 664 -1988 670 1988
rect 704 -1988 710 1988
rect 664 -2000 710 -1988
rect 1122 1988 1168 2000
rect 1122 -1988 1128 1988
rect 1162 -1988 1168 1988
rect 1122 -2000 1168 -1988
rect -1112 -2038 -720 -2032
rect -1112 -2072 -1100 -2038
rect -732 -2072 -720 -2038
rect -1112 -2078 -720 -2072
rect -654 -2038 -262 -2032
rect -654 -2072 -642 -2038
rect -274 -2072 -262 -2038
rect -654 -2078 -262 -2072
rect -196 -2038 196 -2032
rect -196 -2072 -184 -2038
rect 184 -2072 196 -2038
rect -196 -2078 196 -2072
rect 262 -2038 654 -2032
rect 262 -2072 274 -2038
rect 642 -2072 654 -2038
rect 262 -2078 654 -2072
rect 720 -2038 1112 -2032
rect 720 -2072 732 -2038
rect 1100 -2072 1112 -2038
rect 720 -2078 1112 -2072
<< properties >>
string FIXED_BBOX -343 -1157 343 1157
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 10.0 l 2.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
