magic
tech sky130A
magscale 1 2
timestamp 1713056482
<< nwell >>
rect -2225 -2837 2225 2837
<< pmos >>
rect -2029 118 -29 2618
rect 29 118 2029 2618
rect -2029 -2618 -29 -118
rect 29 -2618 2029 -118
<< pdiff >>
rect -2087 2606 -2029 2618
rect -2087 130 -2075 2606
rect -2041 130 -2029 2606
rect -2087 118 -2029 130
rect -29 2606 29 2618
rect -29 130 -17 2606
rect 17 130 29 2606
rect -29 118 29 130
rect 2029 2606 2087 2618
rect 2029 130 2041 2606
rect 2075 130 2087 2606
rect 2029 118 2087 130
rect -2087 -130 -2029 -118
rect -2087 -2606 -2075 -130
rect -2041 -2606 -2029 -130
rect -2087 -2618 -2029 -2606
rect -29 -130 29 -118
rect -29 -2606 -17 -130
rect 17 -2606 29 -130
rect -29 -2618 29 -2606
rect 2029 -130 2087 -118
rect 2029 -2606 2041 -130
rect 2075 -2606 2087 -130
rect 2029 -2618 2087 -2606
<< pdiffc >>
rect -2075 130 -2041 2606
rect -17 130 17 2606
rect 2041 130 2075 2606
rect -2075 -2606 -2041 -130
rect -17 -2606 17 -130
rect 2041 -2606 2075 -130
<< nsubdiff >>
rect -2189 2767 -2093 2801
rect 2093 2767 2189 2801
rect -2189 2705 -2155 2767
rect 2155 2705 2189 2767
rect -2189 -2767 -2155 -2705
rect 2155 -2767 2189 -2705
rect -2189 -2801 -2093 -2767
rect 2093 -2801 2189 -2767
<< nsubdiffcont >>
rect -2093 2767 2093 2801
rect -2189 -2705 -2155 2705
rect 2155 -2705 2189 2705
rect -2093 -2801 2093 -2767
<< poly >>
rect -2029 2699 -29 2715
rect -2029 2665 -2013 2699
rect -45 2665 -29 2699
rect -2029 2618 -29 2665
rect 29 2699 2029 2715
rect 29 2665 45 2699
rect 2013 2665 2029 2699
rect 29 2618 2029 2665
rect -2029 71 -29 118
rect -2029 37 -2013 71
rect -45 37 -29 71
rect -2029 21 -29 37
rect 29 71 2029 118
rect 29 37 45 71
rect 2013 37 2029 71
rect 29 21 2029 37
rect -2029 -37 -29 -21
rect -2029 -71 -2013 -37
rect -45 -71 -29 -37
rect -2029 -118 -29 -71
rect 29 -37 2029 -21
rect 29 -71 45 -37
rect 2013 -71 2029 -37
rect 29 -118 2029 -71
rect -2029 -2665 -29 -2618
rect -2029 -2699 -2013 -2665
rect -45 -2699 -29 -2665
rect -2029 -2715 -29 -2699
rect 29 -2665 2029 -2618
rect 29 -2699 45 -2665
rect 2013 -2699 2029 -2665
rect 29 -2715 2029 -2699
<< polycont >>
rect -2013 2665 -45 2699
rect 45 2665 2013 2699
rect -2013 37 -45 71
rect 45 37 2013 71
rect -2013 -71 -45 -37
rect 45 -71 2013 -37
rect -2013 -2699 -45 -2665
rect 45 -2699 2013 -2665
<< locali >>
rect -2189 2767 -2093 2801
rect 2093 2767 2189 2801
rect -2189 2705 -2155 2767
rect 2155 2705 2189 2767
rect -2029 2665 -2013 2699
rect -45 2665 -29 2699
rect 29 2665 45 2699
rect 2013 2665 2029 2699
rect -2075 2606 -2041 2622
rect -2075 114 -2041 130
rect -17 2606 17 2622
rect -17 114 17 130
rect 2041 2606 2075 2622
rect 2041 114 2075 130
rect -2029 37 -2013 71
rect -45 37 -29 71
rect 29 37 45 71
rect 2013 37 2029 71
rect -2029 -71 -2013 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 2013 -71 2029 -37
rect -2075 -130 -2041 -114
rect -2075 -2622 -2041 -2606
rect -17 -130 17 -114
rect -17 -2622 17 -2606
rect 2041 -130 2075 -114
rect 2041 -2622 2075 -2606
rect -2029 -2699 -2013 -2665
rect -45 -2699 -29 -2665
rect 29 -2699 45 -2665
rect 2013 -2699 2029 -2665
rect -2189 -2767 -2155 -2705
rect 2155 -2767 2189 -2705
rect -2189 -2801 -2093 -2767
rect 2093 -2801 2189 -2767
<< viali >>
rect -2013 2665 -45 2699
rect 45 2665 2013 2699
rect -2075 130 -2041 2606
rect -17 130 17 2606
rect 2041 130 2075 2606
rect -2013 37 -45 71
rect 45 37 2013 71
rect -2013 -71 -45 -37
rect 45 -71 2013 -37
rect -2075 -2606 -2041 -130
rect -17 -2606 17 -130
rect 2041 -2606 2075 -130
rect -2013 -2699 -45 -2665
rect 45 -2699 2013 -2665
<< metal1 >>
rect -2025 2699 -33 2705
rect -2025 2665 -2013 2699
rect -45 2665 -33 2699
rect -2025 2659 -33 2665
rect 33 2699 2025 2705
rect 33 2665 45 2699
rect 2013 2665 2025 2699
rect 33 2659 2025 2665
rect -2081 2606 -2035 2618
rect -2081 130 -2075 2606
rect -2041 130 -2035 2606
rect -2081 118 -2035 130
rect -23 2606 23 2618
rect -23 130 -17 2606
rect 17 130 23 2606
rect -23 118 23 130
rect 2035 2606 2081 2618
rect 2035 130 2041 2606
rect 2075 130 2081 2606
rect 2035 118 2081 130
rect -2025 71 -33 77
rect -2025 37 -2013 71
rect -45 37 -33 71
rect -2025 31 -33 37
rect 33 71 2025 77
rect 33 37 45 71
rect 2013 37 2025 71
rect 33 31 2025 37
rect -2025 -37 -33 -31
rect -2025 -71 -2013 -37
rect -45 -71 -33 -37
rect -2025 -77 -33 -71
rect 33 -37 2025 -31
rect 33 -71 45 -37
rect 2013 -71 2025 -37
rect 33 -77 2025 -71
rect -2081 -130 -2035 -118
rect -2081 -2606 -2075 -130
rect -2041 -2606 -2035 -130
rect -2081 -2618 -2035 -2606
rect -23 -130 23 -118
rect -23 -2606 -17 -130
rect 17 -2606 23 -130
rect -23 -2618 23 -2606
rect 2035 -130 2081 -118
rect 2035 -2606 2041 -130
rect 2075 -2606 2081 -130
rect 2035 -2618 2081 -2606
rect -2025 -2665 -33 -2659
rect -2025 -2699 -2013 -2665
rect -45 -2699 -33 -2665
rect -2025 -2705 -33 -2699
rect 33 -2665 2025 -2659
rect 33 -2699 45 -2665
rect 2013 -2699 2025 -2665
rect 33 -2705 2025 -2699
<< properties >>
string FIXED_BBOX -2172 -2784 2172 2784
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 12.5 l 10.0 m 2 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
