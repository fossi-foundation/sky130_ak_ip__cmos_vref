magic
tech sky130A
magscale 1 2
timestamp 1713046718
<< pwell >>
rect -396 -11191 396 11191
<< nmos >>
rect -200 8981 200 10981
rect -200 6763 200 8763
rect -200 4545 200 6545
rect -200 2327 200 4327
rect -200 109 200 2109
rect -200 -2109 200 -109
rect -200 -4327 200 -2327
rect -200 -6545 200 -4545
rect -200 -8763 200 -6763
rect -200 -10981 200 -8981
<< ndiff >>
rect -258 10969 -200 10981
rect -258 8993 -246 10969
rect -212 8993 -200 10969
rect -258 8981 -200 8993
rect 200 10969 258 10981
rect 200 8993 212 10969
rect 246 8993 258 10969
rect 200 8981 258 8993
rect -258 8751 -200 8763
rect -258 6775 -246 8751
rect -212 6775 -200 8751
rect -258 6763 -200 6775
rect 200 8751 258 8763
rect 200 6775 212 8751
rect 246 6775 258 8751
rect 200 6763 258 6775
rect -258 6533 -200 6545
rect -258 4557 -246 6533
rect -212 4557 -200 6533
rect -258 4545 -200 4557
rect 200 6533 258 6545
rect 200 4557 212 6533
rect 246 4557 258 6533
rect 200 4545 258 4557
rect -258 4315 -200 4327
rect -258 2339 -246 4315
rect -212 2339 -200 4315
rect -258 2327 -200 2339
rect 200 4315 258 4327
rect 200 2339 212 4315
rect 246 2339 258 4315
rect 200 2327 258 2339
rect -258 2097 -200 2109
rect -258 121 -246 2097
rect -212 121 -200 2097
rect -258 109 -200 121
rect 200 2097 258 2109
rect 200 121 212 2097
rect 246 121 258 2097
rect 200 109 258 121
rect -258 -121 -200 -109
rect -258 -2097 -246 -121
rect -212 -2097 -200 -121
rect -258 -2109 -200 -2097
rect 200 -121 258 -109
rect 200 -2097 212 -121
rect 246 -2097 258 -121
rect 200 -2109 258 -2097
rect -258 -2339 -200 -2327
rect -258 -4315 -246 -2339
rect -212 -4315 -200 -2339
rect -258 -4327 -200 -4315
rect 200 -2339 258 -2327
rect 200 -4315 212 -2339
rect 246 -4315 258 -2339
rect 200 -4327 258 -4315
rect -258 -4557 -200 -4545
rect -258 -6533 -246 -4557
rect -212 -6533 -200 -4557
rect -258 -6545 -200 -6533
rect 200 -4557 258 -4545
rect 200 -6533 212 -4557
rect 246 -6533 258 -4557
rect 200 -6545 258 -6533
rect -258 -6775 -200 -6763
rect -258 -8751 -246 -6775
rect -212 -8751 -200 -6775
rect -258 -8763 -200 -8751
rect 200 -6775 258 -6763
rect 200 -8751 212 -6775
rect 246 -8751 258 -6775
rect 200 -8763 258 -8751
rect -258 -8993 -200 -8981
rect -258 -10969 -246 -8993
rect -212 -10969 -200 -8993
rect -258 -10981 -200 -10969
rect 200 -8993 258 -8981
rect 200 -10969 212 -8993
rect 246 -10969 258 -8993
rect 200 -10981 258 -10969
<< ndiffc >>
rect -246 8993 -212 10969
rect 212 8993 246 10969
rect -246 6775 -212 8751
rect 212 6775 246 8751
rect -246 4557 -212 6533
rect 212 4557 246 6533
rect -246 2339 -212 4315
rect 212 2339 246 4315
rect -246 121 -212 2097
rect 212 121 246 2097
rect -246 -2097 -212 -121
rect 212 -2097 246 -121
rect -246 -4315 -212 -2339
rect 212 -4315 246 -2339
rect -246 -6533 -212 -4557
rect 212 -6533 246 -4557
rect -246 -8751 -212 -6775
rect 212 -8751 246 -6775
rect -246 -10969 -212 -8993
rect 212 -10969 246 -8993
<< psubdiff >>
rect -360 11121 -264 11155
rect 264 11121 360 11155
rect -360 11059 -326 11121
rect 326 11059 360 11121
rect -360 -11121 -326 -11059
rect 326 -11121 360 -11059
rect -360 -11155 -264 -11121
rect 264 -11155 360 -11121
<< psubdiffcont >>
rect -264 11121 264 11155
rect -360 -11059 -326 11059
rect 326 -11059 360 11059
rect -264 -11155 264 -11121
<< poly >>
rect -200 11053 200 11069
rect -200 11019 -184 11053
rect 184 11019 200 11053
rect -200 10981 200 11019
rect -200 8943 200 8981
rect -200 8909 -184 8943
rect 184 8909 200 8943
rect -200 8893 200 8909
rect -200 8835 200 8851
rect -200 8801 -184 8835
rect 184 8801 200 8835
rect -200 8763 200 8801
rect -200 6725 200 6763
rect -200 6691 -184 6725
rect 184 6691 200 6725
rect -200 6675 200 6691
rect -200 6617 200 6633
rect -200 6583 -184 6617
rect 184 6583 200 6617
rect -200 6545 200 6583
rect -200 4507 200 4545
rect -200 4473 -184 4507
rect 184 4473 200 4507
rect -200 4457 200 4473
rect -200 4399 200 4415
rect -200 4365 -184 4399
rect 184 4365 200 4399
rect -200 4327 200 4365
rect -200 2289 200 2327
rect -200 2255 -184 2289
rect 184 2255 200 2289
rect -200 2239 200 2255
rect -200 2181 200 2197
rect -200 2147 -184 2181
rect 184 2147 200 2181
rect -200 2109 200 2147
rect -200 71 200 109
rect -200 37 -184 71
rect 184 37 200 71
rect -200 21 200 37
rect -200 -37 200 -21
rect -200 -71 -184 -37
rect 184 -71 200 -37
rect -200 -109 200 -71
rect -200 -2147 200 -2109
rect -200 -2181 -184 -2147
rect 184 -2181 200 -2147
rect -200 -2197 200 -2181
rect -200 -2255 200 -2239
rect -200 -2289 -184 -2255
rect 184 -2289 200 -2255
rect -200 -2327 200 -2289
rect -200 -4365 200 -4327
rect -200 -4399 -184 -4365
rect 184 -4399 200 -4365
rect -200 -4415 200 -4399
rect -200 -4473 200 -4457
rect -200 -4507 -184 -4473
rect 184 -4507 200 -4473
rect -200 -4545 200 -4507
rect -200 -6583 200 -6545
rect -200 -6617 -184 -6583
rect 184 -6617 200 -6583
rect -200 -6633 200 -6617
rect -200 -6691 200 -6675
rect -200 -6725 -184 -6691
rect 184 -6725 200 -6691
rect -200 -6763 200 -6725
rect -200 -8801 200 -8763
rect -200 -8835 -184 -8801
rect 184 -8835 200 -8801
rect -200 -8851 200 -8835
rect -200 -8909 200 -8893
rect -200 -8943 -184 -8909
rect 184 -8943 200 -8909
rect -200 -8981 200 -8943
rect -200 -11019 200 -10981
rect -200 -11053 -184 -11019
rect 184 -11053 200 -11019
rect -200 -11069 200 -11053
<< polycont >>
rect -184 11019 184 11053
rect -184 8909 184 8943
rect -184 8801 184 8835
rect -184 6691 184 6725
rect -184 6583 184 6617
rect -184 4473 184 4507
rect -184 4365 184 4399
rect -184 2255 184 2289
rect -184 2147 184 2181
rect -184 37 184 71
rect -184 -71 184 -37
rect -184 -2181 184 -2147
rect -184 -2289 184 -2255
rect -184 -4399 184 -4365
rect -184 -4507 184 -4473
rect -184 -6617 184 -6583
rect -184 -6725 184 -6691
rect -184 -8835 184 -8801
rect -184 -8943 184 -8909
rect -184 -11053 184 -11019
<< locali >>
rect -360 11121 -264 11155
rect 264 11121 360 11155
rect -360 11059 -326 11121
rect 326 11059 360 11121
rect -200 11019 -184 11053
rect 184 11019 200 11053
rect -246 10969 -212 10985
rect -246 8977 -212 8993
rect 212 10969 246 10985
rect 212 8977 246 8993
rect -200 8909 -184 8943
rect 184 8909 200 8943
rect -200 8801 -184 8835
rect 184 8801 200 8835
rect -246 8751 -212 8767
rect -246 6759 -212 6775
rect 212 8751 246 8767
rect 212 6759 246 6775
rect -200 6691 -184 6725
rect 184 6691 200 6725
rect -200 6583 -184 6617
rect 184 6583 200 6617
rect -246 6533 -212 6549
rect -246 4541 -212 4557
rect 212 6533 246 6549
rect 212 4541 246 4557
rect -200 4473 -184 4507
rect 184 4473 200 4507
rect -200 4365 -184 4399
rect 184 4365 200 4399
rect -246 4315 -212 4331
rect -246 2323 -212 2339
rect 212 4315 246 4331
rect 212 2323 246 2339
rect -200 2255 -184 2289
rect 184 2255 200 2289
rect -200 2147 -184 2181
rect 184 2147 200 2181
rect -246 2097 -212 2113
rect -246 105 -212 121
rect 212 2097 246 2113
rect 212 105 246 121
rect -200 37 -184 71
rect 184 37 200 71
rect -200 -71 -184 -37
rect 184 -71 200 -37
rect -246 -121 -212 -105
rect -246 -2113 -212 -2097
rect 212 -121 246 -105
rect 212 -2113 246 -2097
rect -200 -2181 -184 -2147
rect 184 -2181 200 -2147
rect -200 -2289 -184 -2255
rect 184 -2289 200 -2255
rect -246 -2339 -212 -2323
rect -246 -4331 -212 -4315
rect 212 -2339 246 -2323
rect 212 -4331 246 -4315
rect -200 -4399 -184 -4365
rect 184 -4399 200 -4365
rect -200 -4507 -184 -4473
rect 184 -4507 200 -4473
rect -246 -4557 -212 -4541
rect -246 -6549 -212 -6533
rect 212 -4557 246 -4541
rect 212 -6549 246 -6533
rect -200 -6617 -184 -6583
rect 184 -6617 200 -6583
rect -200 -6725 -184 -6691
rect 184 -6725 200 -6691
rect -246 -6775 -212 -6759
rect -246 -8767 -212 -8751
rect 212 -6775 246 -6759
rect 212 -8767 246 -8751
rect -200 -8835 -184 -8801
rect 184 -8835 200 -8801
rect -200 -8943 -184 -8909
rect 184 -8943 200 -8909
rect -246 -8993 -212 -8977
rect -246 -10985 -212 -10969
rect 212 -8993 246 -8977
rect 212 -10985 246 -10969
rect -200 -11053 -184 -11019
rect 184 -11053 200 -11019
rect -360 -11121 -326 -11059
rect 326 -11121 360 -11059
rect -360 -11155 -264 -11121
rect 264 -11155 360 -11121
<< viali >>
rect -184 11019 184 11053
rect -246 8993 -212 10969
rect 212 8993 246 10969
rect -184 8909 184 8943
rect -184 8801 184 8835
rect -246 6775 -212 8751
rect 212 6775 246 8751
rect -184 6691 184 6725
rect -184 6583 184 6617
rect -246 4557 -212 6533
rect 212 4557 246 6533
rect -184 4473 184 4507
rect -184 4365 184 4399
rect -246 2339 -212 4315
rect 212 2339 246 4315
rect -184 2255 184 2289
rect -184 2147 184 2181
rect -246 121 -212 2097
rect 212 121 246 2097
rect -184 37 184 71
rect -184 -71 184 -37
rect -246 -2097 -212 -121
rect 212 -2097 246 -121
rect -184 -2181 184 -2147
rect -184 -2289 184 -2255
rect -246 -4315 -212 -2339
rect 212 -4315 246 -2339
rect -184 -4399 184 -4365
rect -184 -4507 184 -4473
rect -246 -6533 -212 -4557
rect 212 -6533 246 -4557
rect -184 -6617 184 -6583
rect -184 -6725 184 -6691
rect -246 -8751 -212 -6775
rect 212 -8751 246 -6775
rect -184 -8835 184 -8801
rect -184 -8943 184 -8909
rect -246 -10969 -212 -8993
rect 212 -10969 246 -8993
rect -184 -11053 184 -11019
<< metal1 >>
rect -196 11053 196 11059
rect -196 11019 -184 11053
rect 184 11019 196 11053
rect -196 11013 196 11019
rect -252 10969 -206 10981
rect -252 8993 -246 10969
rect -212 8993 -206 10969
rect -252 8981 -206 8993
rect 206 10969 252 10981
rect 206 8993 212 10969
rect 246 8993 252 10969
rect 206 8981 252 8993
rect -196 8943 196 8949
rect -196 8909 -184 8943
rect 184 8909 196 8943
rect -196 8903 196 8909
rect -196 8835 196 8841
rect -196 8801 -184 8835
rect 184 8801 196 8835
rect -196 8795 196 8801
rect -252 8751 -206 8763
rect -252 6775 -246 8751
rect -212 6775 -206 8751
rect -252 6763 -206 6775
rect 206 8751 252 8763
rect 206 6775 212 8751
rect 246 6775 252 8751
rect 206 6763 252 6775
rect -196 6725 196 6731
rect -196 6691 -184 6725
rect 184 6691 196 6725
rect -196 6685 196 6691
rect -196 6617 196 6623
rect -196 6583 -184 6617
rect 184 6583 196 6617
rect -196 6577 196 6583
rect -252 6533 -206 6545
rect -252 4557 -246 6533
rect -212 4557 -206 6533
rect -252 4545 -206 4557
rect 206 6533 252 6545
rect 206 4557 212 6533
rect 246 4557 252 6533
rect 206 4545 252 4557
rect -196 4507 196 4513
rect -196 4473 -184 4507
rect 184 4473 196 4507
rect -196 4467 196 4473
rect -196 4399 196 4405
rect -196 4365 -184 4399
rect 184 4365 196 4399
rect -196 4359 196 4365
rect -252 4315 -206 4327
rect -252 2339 -246 4315
rect -212 2339 -206 4315
rect -252 2327 -206 2339
rect 206 4315 252 4327
rect 206 2339 212 4315
rect 246 2339 252 4315
rect 206 2327 252 2339
rect -196 2289 196 2295
rect -196 2255 -184 2289
rect 184 2255 196 2289
rect -196 2249 196 2255
rect -196 2181 196 2187
rect -196 2147 -184 2181
rect 184 2147 196 2181
rect -196 2141 196 2147
rect -252 2097 -206 2109
rect -252 121 -246 2097
rect -212 121 -206 2097
rect -252 109 -206 121
rect 206 2097 252 2109
rect 206 121 212 2097
rect 246 121 252 2097
rect 206 109 252 121
rect -196 71 196 77
rect -196 37 -184 71
rect 184 37 196 71
rect -196 31 196 37
rect -196 -37 196 -31
rect -196 -71 -184 -37
rect 184 -71 196 -37
rect -196 -77 196 -71
rect -252 -121 -206 -109
rect -252 -2097 -246 -121
rect -212 -2097 -206 -121
rect -252 -2109 -206 -2097
rect 206 -121 252 -109
rect 206 -2097 212 -121
rect 246 -2097 252 -121
rect 206 -2109 252 -2097
rect -196 -2147 196 -2141
rect -196 -2181 -184 -2147
rect 184 -2181 196 -2147
rect -196 -2187 196 -2181
rect -196 -2255 196 -2249
rect -196 -2289 -184 -2255
rect 184 -2289 196 -2255
rect -196 -2295 196 -2289
rect -252 -2339 -206 -2327
rect -252 -4315 -246 -2339
rect -212 -4315 -206 -2339
rect -252 -4327 -206 -4315
rect 206 -2339 252 -2327
rect 206 -4315 212 -2339
rect 246 -4315 252 -2339
rect 206 -4327 252 -4315
rect -196 -4365 196 -4359
rect -196 -4399 -184 -4365
rect 184 -4399 196 -4365
rect -196 -4405 196 -4399
rect -196 -4473 196 -4467
rect -196 -4507 -184 -4473
rect 184 -4507 196 -4473
rect -196 -4513 196 -4507
rect -252 -4557 -206 -4545
rect -252 -6533 -246 -4557
rect -212 -6533 -206 -4557
rect -252 -6545 -206 -6533
rect 206 -4557 252 -4545
rect 206 -6533 212 -4557
rect 246 -6533 252 -4557
rect 206 -6545 252 -6533
rect -196 -6583 196 -6577
rect -196 -6617 -184 -6583
rect 184 -6617 196 -6583
rect -196 -6623 196 -6617
rect -196 -6691 196 -6685
rect -196 -6725 -184 -6691
rect 184 -6725 196 -6691
rect -196 -6731 196 -6725
rect -252 -6775 -206 -6763
rect -252 -8751 -246 -6775
rect -212 -8751 -206 -6775
rect -252 -8763 -206 -8751
rect 206 -6775 252 -6763
rect 206 -8751 212 -6775
rect 246 -8751 252 -6775
rect 206 -8763 252 -8751
rect -196 -8801 196 -8795
rect -196 -8835 -184 -8801
rect 184 -8835 196 -8801
rect -196 -8841 196 -8835
rect -196 -8909 196 -8903
rect -196 -8943 -184 -8909
rect 184 -8943 196 -8909
rect -196 -8949 196 -8943
rect -252 -8993 -206 -8981
rect -252 -10969 -246 -8993
rect -212 -10969 -206 -8993
rect -252 -10981 -206 -10969
rect 206 -8993 252 -8981
rect 206 -10969 212 -8993
rect 246 -10969 252 -8993
rect 206 -10981 252 -10969
rect -196 -11019 196 -11013
rect -196 -11053 -184 -11019
rect 184 -11053 196 -11019
rect -196 -11059 196 -11053
<< properties >>
string FIXED_BBOX -343 -11138 343 11138
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 10.0 l 2.0 m 10 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
