magic
tech sky130A
magscale 1 2
timestamp 1713051387
<< pwell >>
rect -352 -927 352 927
<< psubdiff >>
rect -316 857 -220 891
rect 220 857 316 891
rect -316 795 -282 857
rect 282 795 316 857
rect -316 -857 -282 -795
rect 282 -857 316 -795
rect -316 -891 -220 -857
rect 220 -891 316 -857
<< psubdiffcont >>
rect -220 857 220 891
rect -316 -795 -282 795
rect 282 -795 316 795
rect -220 -891 220 -857
<< xpolycontact >>
rect -186 329 -48 761
rect -186 -761 -48 -329
rect 48 329 186 761
rect 48 -761 186 -329
<< xpolyres >>
rect -186 -329 -48 329
rect 48 -329 186 329
<< locali >>
rect -316 857 -220 891
rect 220 857 316 891
rect -316 795 -282 857
rect 282 795 316 857
rect -316 -857 -282 -795
rect 282 -857 316 -795
rect -316 -891 -220 -857
rect 220 -891 316 -857
<< viali >>
rect -170 346 -64 743
rect 64 346 170 743
rect -170 -743 -64 -346
rect 64 -743 170 -346
<< metal1 >>
rect -176 743 -58 755
rect -176 346 -170 743
rect -64 346 -58 743
rect -176 334 -58 346
rect 58 743 176 755
rect 58 346 64 743
rect 170 346 176 743
rect 58 334 176 346
rect -176 -346 -58 -334
rect -176 -743 -170 -346
rect -64 -743 -58 -346
rect -176 -755 -58 -743
rect 58 -346 176 -334
rect 58 -743 64 -346
rect 170 -743 176 -346
rect 58 -755 176 -743
<< properties >>
string FIXED_BBOX -299 -874 299 874
string gencell sky130_fd_pr__res_xhigh_po_0p69
string library sky130
string parameters w 0.69 l 3.45 m 1 nx 2 wmin 0.690 lmin 0.50 rho 2000 val 10.545k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.690 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
