magic
tech sky130A
magscale 1 2
timestamp 1713212409
<< pwell >>
rect -1999 -1460 1999 1460
<< nmos >>
rect -1803 -1250 -1403 1250
rect -1345 -1250 -945 1250
rect -887 -1250 -487 1250
rect -429 -1250 -29 1250
rect 29 -1250 429 1250
rect 487 -1250 887 1250
rect 945 -1250 1345 1250
rect 1403 -1250 1803 1250
<< ndiff >>
rect -1861 1238 -1803 1250
rect -1861 -1238 -1849 1238
rect -1815 -1238 -1803 1238
rect -1861 -1250 -1803 -1238
rect -1403 1238 -1345 1250
rect -1403 -1238 -1391 1238
rect -1357 -1238 -1345 1238
rect -1403 -1250 -1345 -1238
rect -945 1238 -887 1250
rect -945 -1238 -933 1238
rect -899 -1238 -887 1238
rect -945 -1250 -887 -1238
rect -487 1238 -429 1250
rect -487 -1238 -475 1238
rect -441 -1238 -429 1238
rect -487 -1250 -429 -1238
rect -29 1238 29 1250
rect -29 -1238 -17 1238
rect 17 -1238 29 1238
rect -29 -1250 29 -1238
rect 429 1238 487 1250
rect 429 -1238 441 1238
rect 475 -1238 487 1238
rect 429 -1250 487 -1238
rect 887 1238 945 1250
rect 887 -1238 899 1238
rect 933 -1238 945 1238
rect 887 -1250 945 -1238
rect 1345 1238 1403 1250
rect 1345 -1238 1357 1238
rect 1391 -1238 1403 1238
rect 1345 -1250 1403 -1238
rect 1803 1238 1861 1250
rect 1803 -1238 1815 1238
rect 1849 -1238 1861 1238
rect 1803 -1250 1861 -1238
<< ndiffc >>
rect -1849 -1238 -1815 1238
rect -1391 -1238 -1357 1238
rect -933 -1238 -899 1238
rect -475 -1238 -441 1238
rect -17 -1238 17 1238
rect 441 -1238 475 1238
rect 899 -1238 933 1238
rect 1357 -1238 1391 1238
rect 1815 -1238 1849 1238
<< psubdiff >>
rect -1963 1390 -1867 1424
rect 1867 1390 1963 1424
rect -1963 1328 -1929 1390
rect 1929 1328 1963 1390
rect -1963 -1390 -1929 -1328
rect 1929 -1390 1963 -1328
rect -1963 -1424 -1867 -1390
rect 1867 -1424 1963 -1390
<< psubdiffcont >>
rect -1867 1390 1867 1424
rect -1963 -1328 -1929 1328
rect 1929 -1328 1963 1328
rect -1867 -1424 1867 -1390
<< poly >>
rect -1803 1322 -1403 1338
rect -1803 1288 -1787 1322
rect -1419 1288 -1403 1322
rect -1803 1250 -1403 1288
rect -1345 1322 -945 1338
rect -1345 1288 -1329 1322
rect -961 1288 -945 1322
rect -1345 1250 -945 1288
rect -887 1322 -487 1338
rect -887 1288 -871 1322
rect -503 1288 -487 1322
rect -887 1250 -487 1288
rect -429 1322 -29 1338
rect -429 1288 -413 1322
rect -45 1288 -29 1322
rect -429 1250 -29 1288
rect 29 1322 429 1338
rect 29 1288 45 1322
rect 413 1288 429 1322
rect 29 1250 429 1288
rect 487 1322 887 1338
rect 487 1288 503 1322
rect 871 1288 887 1322
rect 487 1250 887 1288
rect 945 1322 1345 1338
rect 945 1288 961 1322
rect 1329 1288 1345 1322
rect 945 1250 1345 1288
rect 1403 1322 1803 1338
rect 1403 1288 1419 1322
rect 1787 1288 1803 1322
rect 1403 1250 1803 1288
rect -1803 -1288 -1403 -1250
rect -1803 -1322 -1787 -1288
rect -1419 -1322 -1403 -1288
rect -1803 -1338 -1403 -1322
rect -1345 -1288 -945 -1250
rect -1345 -1322 -1329 -1288
rect -961 -1322 -945 -1288
rect -1345 -1338 -945 -1322
rect -887 -1288 -487 -1250
rect -887 -1322 -871 -1288
rect -503 -1322 -487 -1288
rect -887 -1338 -487 -1322
rect -429 -1288 -29 -1250
rect -429 -1322 -413 -1288
rect -45 -1322 -29 -1288
rect -429 -1338 -29 -1322
rect 29 -1288 429 -1250
rect 29 -1322 45 -1288
rect 413 -1322 429 -1288
rect 29 -1338 429 -1322
rect 487 -1288 887 -1250
rect 487 -1322 503 -1288
rect 871 -1322 887 -1288
rect 487 -1338 887 -1322
rect 945 -1288 1345 -1250
rect 945 -1322 961 -1288
rect 1329 -1322 1345 -1288
rect 945 -1338 1345 -1322
rect 1403 -1288 1803 -1250
rect 1403 -1322 1419 -1288
rect 1787 -1322 1803 -1288
rect 1403 -1338 1803 -1322
<< polycont >>
rect -1787 1288 -1419 1322
rect -1329 1288 -961 1322
rect -871 1288 -503 1322
rect -413 1288 -45 1322
rect 45 1288 413 1322
rect 503 1288 871 1322
rect 961 1288 1329 1322
rect 1419 1288 1787 1322
rect -1787 -1322 -1419 -1288
rect -1329 -1322 -961 -1288
rect -871 -1322 -503 -1288
rect -413 -1322 -45 -1288
rect 45 -1322 413 -1288
rect 503 -1322 871 -1288
rect 961 -1322 1329 -1288
rect 1419 -1322 1787 -1288
<< locali >>
rect -1963 1390 -1867 1424
rect 1867 1390 1963 1424
rect -1963 1328 -1929 1390
rect 1929 1328 1963 1390
rect -1803 1288 -1787 1322
rect -1419 1288 -1403 1322
rect -1345 1288 -1329 1322
rect -961 1288 -945 1322
rect -887 1288 -871 1322
rect -503 1288 -487 1322
rect -429 1288 -413 1322
rect -45 1288 -29 1322
rect 29 1288 45 1322
rect 413 1288 429 1322
rect 487 1288 503 1322
rect 871 1288 887 1322
rect 945 1288 961 1322
rect 1329 1288 1345 1322
rect 1403 1288 1419 1322
rect 1787 1288 1803 1322
rect -1849 1238 -1815 1254
rect -1849 -1254 -1815 -1238
rect -1391 1238 -1357 1254
rect -1391 -1254 -1357 -1238
rect -933 1238 -899 1254
rect -933 -1254 -899 -1238
rect -475 1238 -441 1254
rect -475 -1254 -441 -1238
rect -17 1238 17 1254
rect -17 -1254 17 -1238
rect 441 1238 475 1254
rect 441 -1254 475 -1238
rect 899 1238 933 1254
rect 899 -1254 933 -1238
rect 1357 1238 1391 1254
rect 1357 -1254 1391 -1238
rect 1815 1238 1849 1254
rect 1815 -1254 1849 -1238
rect -1803 -1322 -1787 -1288
rect -1419 -1322 -1403 -1288
rect -1345 -1322 -1329 -1288
rect -961 -1322 -945 -1288
rect -887 -1322 -871 -1288
rect -503 -1322 -487 -1288
rect -429 -1322 -413 -1288
rect -45 -1322 -29 -1288
rect 29 -1322 45 -1288
rect 413 -1322 429 -1288
rect 487 -1322 503 -1288
rect 871 -1322 887 -1288
rect 945 -1322 961 -1288
rect 1329 -1322 1345 -1288
rect 1403 -1322 1419 -1288
rect 1787 -1322 1803 -1288
rect -1963 -1390 -1929 -1328
rect 1929 -1390 1963 -1328
rect -1963 -1424 -1867 -1390
rect 1867 -1424 1963 -1390
<< viali >>
rect -1787 1288 -1419 1322
rect -1329 1288 -961 1322
rect -871 1288 -503 1322
rect -413 1288 -45 1322
rect 45 1288 413 1322
rect 503 1288 871 1322
rect 961 1288 1329 1322
rect 1419 1288 1787 1322
rect -1849 -1238 -1815 1238
rect -1391 -1238 -1357 1238
rect -933 -1238 -899 1238
rect -475 -1238 -441 1238
rect -17 -1238 17 1238
rect 441 -1238 475 1238
rect 899 -1238 933 1238
rect 1357 -1238 1391 1238
rect 1815 -1238 1849 1238
rect -1787 -1322 -1419 -1288
rect -1329 -1322 -961 -1288
rect -871 -1322 -503 -1288
rect -413 -1322 -45 -1288
rect 45 -1322 413 -1288
rect 503 -1322 871 -1288
rect 961 -1322 1329 -1288
rect 1419 -1322 1787 -1288
<< metal1 >>
rect -1799 1322 -1407 1328
rect -1799 1288 -1787 1322
rect -1419 1288 -1407 1322
rect -1799 1282 -1407 1288
rect -1341 1322 -949 1328
rect -1341 1288 -1329 1322
rect -961 1288 -949 1322
rect -1341 1282 -949 1288
rect -883 1322 -491 1328
rect -883 1288 -871 1322
rect -503 1288 -491 1322
rect -883 1282 -491 1288
rect -425 1322 -33 1328
rect -425 1288 -413 1322
rect -45 1288 -33 1322
rect -425 1282 -33 1288
rect 33 1322 425 1328
rect 33 1288 45 1322
rect 413 1288 425 1322
rect 33 1282 425 1288
rect 491 1322 883 1328
rect 491 1288 503 1322
rect 871 1288 883 1322
rect 491 1282 883 1288
rect 949 1322 1341 1328
rect 949 1288 961 1322
rect 1329 1288 1341 1322
rect 949 1282 1341 1288
rect 1407 1322 1799 1328
rect 1407 1288 1419 1322
rect 1787 1288 1799 1322
rect 1407 1282 1799 1288
rect -1855 1238 -1809 1250
rect -1855 -1238 -1849 1238
rect -1815 -1238 -1809 1238
rect -1855 -1250 -1809 -1238
rect -1397 1238 -1351 1250
rect -1397 -1238 -1391 1238
rect -1357 -1238 -1351 1238
rect -1397 -1250 -1351 -1238
rect -939 1238 -893 1250
rect -939 -1238 -933 1238
rect -899 -1238 -893 1238
rect -939 -1250 -893 -1238
rect -481 1238 -435 1250
rect -481 -1238 -475 1238
rect -441 -1238 -435 1238
rect -481 -1250 -435 -1238
rect -23 1238 23 1250
rect -23 -1238 -17 1238
rect 17 -1238 23 1238
rect -23 -1250 23 -1238
rect 435 1238 481 1250
rect 435 -1238 441 1238
rect 475 -1238 481 1238
rect 435 -1250 481 -1238
rect 893 1238 939 1250
rect 893 -1238 899 1238
rect 933 -1238 939 1238
rect 893 -1250 939 -1238
rect 1351 1238 1397 1250
rect 1351 -1238 1357 1238
rect 1391 -1238 1397 1238
rect 1351 -1250 1397 -1238
rect 1809 1238 1855 1250
rect 1809 -1238 1815 1238
rect 1849 -1238 1855 1238
rect 1809 -1250 1855 -1238
rect -1799 -1288 -1407 -1282
rect -1799 -1322 -1787 -1288
rect -1419 -1322 -1407 -1288
rect -1799 -1328 -1407 -1322
rect -1341 -1288 -949 -1282
rect -1341 -1322 -1329 -1288
rect -961 -1322 -949 -1288
rect -1341 -1328 -949 -1322
rect -883 -1288 -491 -1282
rect -883 -1322 -871 -1288
rect -503 -1322 -491 -1288
rect -883 -1328 -491 -1322
rect -425 -1288 -33 -1282
rect -425 -1322 -413 -1288
rect -45 -1322 -33 -1288
rect -425 -1328 -33 -1322
rect 33 -1288 425 -1282
rect 33 -1322 45 -1288
rect 413 -1322 425 -1288
rect 33 -1328 425 -1322
rect 491 -1288 883 -1282
rect 491 -1322 503 -1288
rect 871 -1322 883 -1288
rect 491 -1328 883 -1322
rect 949 -1288 1341 -1282
rect 949 -1322 961 -1288
rect 1329 -1322 1341 -1288
rect 949 -1328 1341 -1322
rect 1407 -1288 1799 -1282
rect 1407 -1322 1419 -1288
rect 1787 -1322 1799 -1288
rect 1407 -1328 1799 -1322
<< properties >>
string FIXED_BBOX -1946 -1407 1946 1407
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 12.5 l 2.0 m 1 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
