magic
tech sky130A
timestamp 1713212409
<< pwell >>
rect -348 -605 348 605
<< nmos >>
rect -250 -500 250 500
<< ndiff >>
rect -279 494 -250 500
rect -279 -494 -273 494
rect -256 -494 -250 494
rect -279 -500 -250 -494
rect 250 494 279 500
rect 250 -494 256 494
rect 273 -494 279 494
rect 250 -500 279 -494
<< ndiffc >>
rect -273 -494 -256 494
rect 256 -494 273 494
<< psubdiff >>
rect -330 570 -282 587
rect 282 570 330 587
rect -330 539 -313 570
rect 313 539 330 570
rect -330 -570 -313 -539
rect 313 -570 330 -539
rect -330 -587 -282 -570
rect 282 -587 330 -570
<< psubdiffcont >>
rect -282 570 282 587
rect -330 -539 -313 539
rect 313 -539 330 539
rect -282 -587 282 -570
<< poly >>
rect -250 536 250 544
rect -250 519 -242 536
rect 242 519 250 536
rect -250 500 250 519
rect -250 -519 250 -500
rect -250 -536 -242 -519
rect 242 -536 250 -519
rect -250 -544 250 -536
<< polycont >>
rect -242 519 242 536
rect -242 -536 242 -519
<< locali >>
rect -330 570 -282 587
rect 282 570 330 587
rect -330 539 -313 570
rect 313 539 330 570
rect -250 519 -242 536
rect 242 519 250 536
rect -273 494 -256 502
rect -273 -502 -256 -494
rect 256 494 273 502
rect 256 -502 273 -494
rect -250 -536 -242 -519
rect 242 -536 250 -519
rect -330 -570 -313 -539
rect 313 -570 330 -539
rect -330 -587 -282 -570
rect 282 -587 330 -570
<< viali >>
rect -242 519 242 536
rect -273 -494 -256 494
rect 256 -494 273 494
rect -242 -536 242 -519
<< metal1 >>
rect -248 536 248 539
rect -248 519 -242 536
rect 242 519 248 536
rect -248 516 248 519
rect -276 494 -253 500
rect -276 -494 -273 494
rect -256 -494 -253 494
rect -276 -500 -253 -494
rect 253 494 276 500
rect 253 -494 256 494
rect 273 -494 276 494
rect 253 -500 276 -494
rect -248 -519 248 -516
rect -248 -536 -242 -519
rect 242 -536 248 -519
rect -248 -539 248 -536
<< properties >>
string FIXED_BBOX -321 -578 321 578
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 10 l 5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
